module C3540 ( G1_0_gat, G13_1_gat, G20_2_gat, G33_3_gat, G41_4_gat, G45_5_gat, G50_6_gat, G58_7_gat, G68_8_gat, G77_9_gat, G87_10_gat, G97_11_gat, G107_12_gat, G116_13_gat, G124_14_gat, G125_15_gat, G128_16_gat, G132_17_gat, G137_18_gat, G143_19_gat, G150_20_gat, G159_21_gat, G169_22_gat, G179_23_gat, G190_24_gat, G200_25_gat, G213_26_gat, G222_27_gat, G223_28_gat, G226_29_gat, G232_30_gat, G238_31_gat, G244_32_gat, G250_33_gat, G257_34_gat, G264_35_gat, G270_36_gat, G274_37_gat, G283_38_gat, G294_39_gat, G303_40_gat, G311_41_gat, G317_42_gat, G322_43_gat, G326_44_gat, G329_45_gat, G330_46_gat, G343_47_gat, G1698_48_gat, G2897_49_gat, G353_405_gat, G355_399_gat, G361_940_gat, G358_1161_gat, G351_1247_gat, G372_1243_gat, G369_1321_gat, G399_1428_gat, G364_1484_gat, G396_1504_gat, G384_1553_gat, G367_1585_gat, G387_1616_gat, G393_1605_gat, G390_1603_gat, G378_1597_gat, G375_1624_gat, G381_1626_gat, G407_1657_gat, G409_1670_gat, G405_1717_gat, G402_1718_gat);

input G1_0_gat;
input G13_1_gat;
input G20_2_gat;
input G33_3_gat;
input G41_4_gat;
input G45_5_gat;
input G50_6_gat;
input G58_7_gat;
input G68_8_gat;
input G77_9_gat;
input G87_10_gat;
input G97_11_gat;
input G107_12_gat;
input G116_13_gat;
input G124_14_gat;
input G125_15_gat;
input G128_16_gat;
input G132_17_gat;
input G137_18_gat;
input G143_19_gat;
input G150_20_gat;
input G159_21_gat;
input G169_22_gat;
input G179_23_gat;
input G190_24_gat;
input G200_25_gat;
input G213_26_gat;
input G222_27_gat;
input G223_28_gat;
input G226_29_gat;
input G232_30_gat;
input G238_31_gat;
input G244_32_gat;
input G250_33_gat;
input G257_34_gat;
input G264_35_gat;
input G270_36_gat;
input G274_37_gat;
input G283_38_gat;
input G294_39_gat;
input G303_40_gat;
input G311_41_gat;
input G317_42_gat;
input G322_43_gat;
input G326_44_gat;
input G329_45_gat;
input G330_46_gat;
input G343_47_gat;
input G1698_48_gat;
input G2897_49_gat;

output G353_405_gat;
output G355_399_gat;
output G361_940_gat;
output G358_1161_gat;
output G351_1247_gat;
output G372_1243_gat;
output G369_1321_gat;
output G399_1428_gat;
output G364_1484_gat;
output G396_1504_gat;
output G384_1553_gat;
output G367_1585_gat;
output G387_1616_gat;
output G393_1605_gat;
output G390_1603_gat;
output G378_1597_gat;
output G375_1624_gat;
output G381_1626_gat;
output G407_1657_gat;
output G409_1670_gat;
output G405_1717_gat;
output G402_1718_gat;

BUFX20 U_g1 (.A(G343_47_gat), .Y(G2868_50_gat) );
BUFX20 U_g2 (.A(G330_46_gat), .Y(G3419_51_gat) );
BUFX20 U_g3 (.A(G270_36_gat), .Y(G2960_52_gat) );
BUFX20 U_g4 (.A(G264_35_gat), .Y(G2957_53_gat) );
AND2XL U_g5 (.A(G264_35_ngat), .B(G257_34_ngat), .Y(G587_54_gat) );
BUFX20 U_g6 (.A(G257_34_gat), .Y(G2950_55_gat) );
BUFX20 U_g7 (.A(G250_33_gat), .Y(G2947_56_gat) );
BUFX20 U_g8 (.A(G244_32_gat), .Y(G2942_57_gat) );
BUFX20 U_g9 (.A(G238_31_gat), .Y(G2939_58_gat) );
BUFX20 U_g10 (.A(G232_30_gat), .Y(G2934_59_gat) );
BUFX20 U_g11 (.A(G226_29_gat), .Y(G2931_60_gat) );
BUFX20 U_g12 (.A(G213_26_gat), .Y(G2865_61_gat) );
BUFX20 U_g13 (.A(G200_25_gat), .Y(G1048_62_gat) );
BUFX20 U_g14 (.A(G190_24_gat), .Y(G1035_63_gat) );
BUFX20 U_g15 (.A(G179_23_gat), .Y(G2478_64_gat) );
BUFX20 U_g16 (.A(G116_13_gat), .Y(G540_65_gat) );
BUFX20 U_g17 (.A(G116_13_gat), .Y(G530_66_gat) );
BUFX20 U_g18 (.A(G107_12_gat), .Y(G907_67_gat) );
BUFX20 U_g19 (.A(G107_12_gat), .Y(G851_68_gat) );
BUFX20 U_g20 (.A(G107_12_gat), .Y(G526_69_gat) );
BUFX20 U_g21 (.A(G107_12_gat), .Y(G517_70_gat) );
BUFX20 U_g22 (.A(G97_11_gat), .Y(G3103_71_gat) );
BUFX20 U_g23 (.A(G97_11_gat), .Y(G3095_72_gat) );
BUFX20 U_g24 (.A(G97_11_gat), .Y(G848_73_gat) );
BUFX20 U_g25 (.A(G97_11_gat), .Y(G845_74_gat) );
BUFX20 U_g26 (.A(G97_11_gat), .Y(G513_75_gat) );
BUFX20 U_g27 (.A(G97_11_gat), .Y(G504_76_gat) );
BUFX20 U_g28 (.A(G87_10_gat), .Y(G842_77_gat) );
BUFX20 U_g29 (.A(G87_10_gat), .Y(G839_78_gat) );
BUFX20 U_g30 (.A(G87_10_gat), .Y(G501_79_gat) );
BUFX20 U_g31 (.A(G87_10_gat), .Y(G492_80_gat) );
BUFX20 U_g32 (.A(G77_9_gat), .Y(G483_81_gat) );
BUFX20 U_g33 (.A(G77_9_gat), .Y(G479_82_gat) );
BUFX20 U_g34 (.A(G77_9_gat), .Y(G476_83_gat) );
BUFX20 U_g35 (.A(G68_8_gat), .Y(G898_84_gat) );
BUFX20 U_g36 (.A(G68_8_gat), .Y(G836_85_gat) );
BUFX20 U_g37 (.A(G68_8_gat), .Y(G833_86_gat) );
BUFX20 U_g38 (.A(G68_8_gat), .Y(G467_87_gat) );
BUFX20 U_g39 (.A(G68_8_gat), .Y(G463_88_gat) );
BUFX20 U_g40 (.A(G68_8_gat), .Y(G460_89_gat) );
BUFX20 U_g41 (.A(G58_7_gat), .Y(G3087_90_gat) );
BUFX20 U_g42 (.A(G58_7_gat), .Y(G3079_91_gat) );
BUFX20 U_g43 (.A(G58_7_gat), .Y(G831_92_gat) );
BUFX20 U_g44 (.A(G58_7_gat), .Y(G828_93_gat) );
BUFX20 U_g45 (.A(G58_7_gat), .Y(G456_94_gat) );
BUFX20 U_g46 (.A(G58_7_gat), .Y(G447_95_gat) );
BUFX20 U_g47 (.A(G50_6_gat), .Y(G826_96_gat) );
BUFX20 U_g48 (.A(G50_6_gat), .Y(G3007_97_gat) );
BUFX20 U_g49 (.A(G50_6_gat), .Y(G442_98_gat) );
BUFX20 U_g50 (.A(G50_6_gat), .Y(G432_99_gat) );
BUFX20 U_g51 (.A(G45_5_gat), .Y(G802_100_gat) );
BUFX20 U_g52 (.A(G45_5_gat), .Y(G799_101_gat) );
AND2XL U_g53 (.A(G45_5_ngat), .B(G41_4_ngat), .Y(G798_102_gat) );
BUFX20 U_g54 (.A(G41_4_gat), .Y(G791_103_gat) );
BUFX20 U_g55 (.A(G33_3_gat), .Y(G2051_104_gat) );
AND2XL U_g56 (.A(G33_3_ngat), .B(G1698_48_ngat), .Y(G1699_105_gat) );
BUFX20 U_g57 (.A(G33_3_gat), .Y(G780_106_gat) );
BUFX20 U_g58 (.A(G33_3_gat), .Y(G776_107_gat) );
BUFX20 U_g59 (.A(G33_3_gat), .Y(G758_108_gat) );
AND2XL U_g60 (.A(G41_4_gat), .B(G33_3_gat), .Y(G788_109_gat) );
BUFX20 U_g61 (.A(G20_2_gat), .Y(G1828_110_gat) );
BUFX20 U_g62 (.A(G20_2_gat), .Y(G1540_111_gat) );
AND2XL U_g63 (.A(G179_23_gat), .B(G20_2_gat), .Y(G1051_112_gat) );
AND2XL U_g64 (.A(G200_25_gat), .B(G20_2_gat), .Y(G1050_113_gat) );
AND2XL U_g65 (.A(G200_25_gat), .B(G20_2_gat), .Y(G1049_114_gat) );
BUFX20 U_g66 (.A(G20_2_gat), .Y(G1032_115_gat) );
BUFX20 U_g67 (.A(G20_2_gat), .Y(G741_116_gat) );
BUFX20 U_g68 (.A(G20_2_gat), .Y(G732_117_gat) );
BUFX20 U_g69 (.A(G20_2_gat), .Y(G736_118_gat) );
BUFX20 U_g70 (.A(G13_1_gat), .Y(G724_119_gat) );
BUFX20 U_g71 (.A(G13_1_gat), .Y(G717_120_gat) );
AND2XL U_g72 (.A(G20_2_gat), .B(G13_1_gat), .Y(G731_121_gat) );
AND3XL U_g73 (.A(G33_3_gat), .B(G20_2_gat), .C(G1_0_gat), .Y(G1827_122_gat) );
AND2XL U_g74 (.A(G13_1_gat), .B(G1_0_gat), .Y(G1826_123_gat) );
BUFX20 U_g75 (.A(G1_0_gat), .Y(G714_124_gat) );
BUFX20 U_g76 (.A(G1_0_gat), .Y(G890_125_gat) );
BUFX20 U_g77 (.A(G1_0_gat), .Y(G704_126_gat) );
BUFX20 U_g78 (.A(G1_0_gat), .Y(G707_127_gat) );
AND2XL U_g79 (.A(G2868_50_ngat), .B(G2865_61_ngat), .Y(G2871_128_gat) );
AND2XL U_g80 (.A(G2868_50_ngat), .B(G2865_61_ngat), .Y(G2874_129_gat) );
BUFX20 U_g81 (.A(G3419_51_gat), .Y(G3425_130_gat) );
BUFX20 U_g82 (.A(G2960_52_gat), .Y(G2964_131_gat) );
AND2XL U_g83 (.A(G530_66_gat), .B(G270_36_gat), .Y(G552_132_gat) );
BUFX20 U_g84 (.A(G2957_53_gat), .Y(G2963_133_gat) );
AND2XL U_g85 (.A(G517_70_gat), .B(G264_35_gat), .Y(G551_134_gat) );
BUFX20 U_g86 (.A(G2950_55_gat), .Y(G2954_135_gat) );
AND2XL U_g87 (.A(G504_76_gat), .B(G257_34_gat), .Y(G550_136_gat) );
AND2XL U_g88 (.A(G587_54_gat), .B(G250_33_gat), .Y(G588_137_gat) );
BUFX20 U_g89 (.A(G2947_56_gat), .Y(G2953_138_gat) );
AND2XL U_g90 (.A(G492_80_gat), .B(G250_33_gat), .Y(G549_139_gat) );
BUFX20 U_g91 (.A(G2942_57_gat), .Y(G2946_140_gat) );
AND2XL U_g92 (.A(G483_81_gat), .B(G244_32_gat), .Y(G548_141_gat) );
BUFX20 U_g93 (.A(G2939_58_gat), .Y(G2945_142_gat) );
AND2XL U_g94 (.A(G467_87_gat), .B(G238_31_gat), .Y(G547_143_gat) );
BUFX20 U_g95 (.A(G2934_59_gat), .Y(G2938_144_gat) );
AND2XL U_g96 (.A(G447_95_gat), .B(G232_30_gat), .Y(G546_145_gat) );
BUFX20 U_g97 (.A(G2931_60_gat), .Y(G2937_146_gat) );
AND2XL U_g98 (.A(G432_99_gat), .B(G226_29_gat), .Y(G545_147_gat) );
AND2XL U_g99 (.A(G1035_63_ngat), .B(G1032_115_ngat), .Y(G1038_148_gat) );
AND2XL U_g100 (.A(G1035_63_ngat), .B(G1032_115_ngat), .Y(G1043_149_gat) );
BUFX20 U_g101 (.A(G2478_64_gat), .Y(G2481_150_gat) );
AND2XL U_g102 (.A(G169_22_ngat), .B(G1540_111_ngat), .Y(G1541_151_gat) );
BUFX20 U_g103 (.A(G540_65_gat), .Y(G3040_152_gat) );
BUFX20 U_g104 (.A(G907_67_gat), .Y(G3098_153_gat) );
BUFX20 U_g105 (.A(G907_67_gat), .Y(G3106_154_gat) );
AND3XL U_g106 (.A(G851_68_gat), .B(G848_73_gat), .C(G842_77_gat), .Y(G905_155_gat) );
AND3XL U_g107 (.A(G851_68_gat), .B(G848_73_gat), .C(G842_77_gat), .Y(G906_156_gat) );
BUFX20 U_g108 (.A(G526_69_gat), .Y(G3037_157_gat) );
AND2XL U_g109 (.A(G526_69_gat), .B(G513_75_gat), .Y(G626_158_gat) );
BUFX20 U_g110 (.A(G3103_71_gat), .Y(G3109_159_gat) );
BUFX20 U_g111 (.A(G3095_72_gat), .Y(G3101_160_gat) );
BUFX20 U_g112 (.A(G513_75_gat), .Y(G3030_161_gat) );
BUFX20 U_g113 (.A(G501_79_gat), .Y(G3027_162_gat) );
BUFX20 U_g114 (.A(G479_82_gat), .Y(G3020_163_gat) );
AND2XL U_g115 (.A(G476_83_gat), .B(G460_89_gat), .Y(G635_164_gat) );
BUFX20 U_g116 (.A(G898_84_gat), .Y(G3082_165_gat) );
BUFX20 U_g117 (.A(G898_84_gat), .Y(G3090_166_gat) );
AND3XL U_g118 (.A(G836_85_gat), .B(G831_92_gat), .C(G826_96_gat), .Y(G625_167_gat) );
AND3XL U_g119 (.A(G836_85_gat), .B(G831_92_gat), .C(G826_96_gat), .Y(G897_168_gat) );
BUFX20 U_g120 (.A(G463_88_gat), .Y(G3017_169_gat) );
AND2XL U_g121 (.A(G463_88_gat), .B(G456_94_gat), .Y(G621_170_gat) );
BUFX20 U_g122 (.A(G3087_90_gat), .Y(G3093_171_gat) );
BUFX20 U_g123 (.A(G3079_91_gat), .Y(G3085_172_gat) );
BUFX20 U_g124 (.A(G456_94_gat), .Y(G3010_173_gat) );
BUFX20 U_g125 (.A(G3007_97_gat), .Y(G3013_174_gat) );
BUFX20 U_g126 (.A(G442_98_gat), .Y(G636_175_gat) );
AND3XL U_g127 (.A(G45_5_gat), .B(G732_117_gat), .C(G717_120_gat), .Y(G896_176_gat) );
BUFX20 U_g128 (.A(G802_100_gat), .Y(G657_177_gat) );
BUFX20 U_g129 (.A(G802_100_gat), .Y(G675_178_gat) );
AND3XL U_g130 (.A(G791_103_gat), .B(G799_101_gat), .C(G714_124_gat), .Y(G816_179_gat) );
AND2XL U_g131 (.A(G799_101_gat), .B(G704_126_gat), .Y(G823_180_gat) );
AND2XL U_g132 (.A(G798_102_gat), .B(G714_124_gat), .Y(G807_181_gat) );
BUFX20 U_g133 (.A(G791_103_gat), .Y(G794_182_gat) );
BUFX20 U_g134 (.A(G1699_105_gat), .Y(G1717_183_gat) );
BUFX20 U_g135 (.A(G1699_105_gat), .Y(G1724_184_gat) );
BUFX20 U_g136 (.A(G1699_105_gat), .Y(G1731_185_gat) );
BUFX20 U_g137 (.A(G1699_105_gat), .Y(G1738_186_gat) );
BUFX20 U_g138 (.A(G1699_105_gat), .Y(G1745_187_gat) );
BUFX20 U_g139 (.A(G1699_105_gat), .Y(G1752_188_gat) );
BUFX20 U_g140 (.A(G1699_105_gat), .Y(G1759_189_gat) );
BUFX20 U_g141 (.A(G1699_105_gat), .Y(G1766_190_gat) );
BUFX20 U_g142 (.A(G780_106_gat), .Y(G784_191_gat) );
BUFX20 U_g143 (.A(G780_106_gat), .Y(G1681_192_gat) );
BUFX20 U_g144 (.A(G776_107_gat), .Y(G1512_193_gat) );
BUFX20 U_g145 (.A(G788_109_gat), .Y(G1790_194_gat) );
BUFX20 U_g146 (.A(G788_109_gat), .Y(G1808_195_gat) );
BUFX20 U_g147 (.A(G1051_112_gat), .Y(G1054_196_gat) );
BUFX20 U_g148 (.A(G1051_112_gat), .Y(G1057_197_gat) );
AND2XL U_g149 (.A(G20_2_ngat), .B(G758_108_ngat), .Y(G759_198_gat) );
BUFX20 U_g150 (.A(G741_116_gat), .Y(G973_199_gat) );
BUFX20 U_g151 (.A(G741_116_gat), .Y(G980_200_gat) );
BUFX20 U_g152 (.A(G741_116_gat), .Y(G987_201_gat) );
BUFX20 U_g153 (.A(G741_116_gat), .Y(G994_202_gat) );
BUFX20 U_g154 (.A(G741_116_gat), .Y(G1001_203_gat) );
BUFX20 U_g155 (.A(G741_116_gat), .Y(G1008_204_gat) );
BUFX20 U_g156 (.A(G741_116_gat), .Y(G1015_205_gat) );
BUFX20 U_g157 (.A(G741_116_gat), .Y(G1022_206_gat) );
AND3XL U_g158 (.A(G732_117_gat), .B(G717_120_gat), .C(G704_126_gat), .Y(G2278_207_gat) );
AND3XL U_g159 (.A(G736_118_gat), .B(G724_119_gat), .C(G707_127_gat), .Y(G860_208_gat) );
AND3XL U_g160 (.A(G736_118_gat), .B(G724_119_gat), .C(G707_127_gat), .Y(G861_209_gat) );
AND2XL U_g161 (.A(G724_119_gat), .B(G707_127_gat), .Y(G864_210_gat) );
BUFX20 U_g162 (.A(G717_120_gat), .Y(G721_211_gat) );
BUFX20 U_g163 (.A(G731_121_gat), .Y(G1772_212_gat) );
AND2XL U_g164 (.A(G1_0_ngat), .B(G2051_104_ngat), .Y(G2052_213_gat) );
AND2XL U_g165 (.A(G1_0_ngat), .B(G1828_110_ngat), .Y(G1829_214_gat) );
AND2XL U_g166 (.A(G1827_122_gat), .B(G1826_123_gat), .Y(G1834_215_gat) );
BUFX20 U_g167 (.A(G890_125_gat), .Y(G893_216_gat) );
BUFX20 U_g168 (.A(G2874_129_gat), .Y(G2877_217_gat) );
AND2XL U_g169 (.A(G2963_133_gat), .B(G2960_52_gat), .Y(G2965_218_gat) );
AND4XL U_g170 (.A(G552_132_gat), .B(G551_134_gat), .C(G550_136_gat), .D(G549_139_gat), .Y(G554_219_gat) );
AND2XL U_g171 (.A(G2964_131_gat), .B(G2957_53_gat), .Y(G2966_220_gat) );
AND2XL U_g172 (.A(G1766_190_gat), .B(G257_34_gat), .Y(G1769_221_gat) );
AND2XL U_g173 (.A(G2953_138_gat), .B(G2950_55_gat), .Y(G2955_222_gat) );
AND2XL U_g174 (.A(G1759_189_gat), .B(G250_33_gat), .Y(G1762_223_gat) );
AND2XL U_g175 (.A(G2954_135_gat), .B(G2947_56_gat), .Y(G2956_224_gat) );
AND2XL U_g176 (.A(G1752_188_gat), .B(G244_32_gat), .Y(G1755_225_gat) );
AND2XL U_g177 (.A(G2945_142_gat), .B(G2942_57_gat), .Y(G560_226_gat) );
AND4XL U_g178 (.A(G548_141_gat), .B(G547_143_gat), .C(G546_145_gat), .D(G545_147_gat), .Y(G553_227_gat) );
AND2XL U_g179 (.A(G1745_187_gat), .B(G238_31_gat), .Y(G1748_228_gat) );
AND2XL U_g180 (.A(G2946_140_gat), .B(G2939_58_gat), .Y(G561_229_gat) );
AND2XL U_g181 (.A(G1738_186_gat), .B(G232_30_gat), .Y(G1741_230_gat) );
AND2XL U_g182 (.A(G2937_146_gat), .B(G2934_59_gat), .Y(G555_231_gat) );
AND2XL U_g183 (.A(G1731_185_gat), .B(G226_29_gat), .Y(G1734_232_gat) );
AND2XL U_g184 (.A(G2938_144_gat), .B(G2931_60_gat), .Y(G556_233_gat) );
AND2XL U_g185 (.A(G1724_184_gat), .B(G223_28_gat), .Y(G1727_234_gat) );
AND2XL U_g186 (.A(G1717_183_gat), .B(G222_27_gat), .Y(G1720_235_gat) );
AND3XL U_g187 (.A(G343_47_gat), .B(G213_26_gat), .C(G2278_207_gat), .Y(G2302_236_gat) );
AND3XL U_g188 (.A(G343_47_gat), .B(G213_26_gat), .C(G2278_207_gat), .Y(G2298_237_gat) );
AND3XL U_g189 (.A(G343_47_gat), .B(G213_26_gat), .C(G2278_207_gat), .Y(G2293_238_gat) );
AND3XL U_g190 (.A(G343_47_gat), .B(G213_26_gat), .C(G2278_207_gat), .Y(G2289_239_gat) );
AND2XL U_g191 (.A(G213_26_gat), .B(G2278_207_gat), .Y(G2288_240_gat) );
AND2XL U_g192 (.A(G213_26_gat), .B(G2278_207_gat), .Y(G2285_241_gat) );
AND2XL U_g193 (.A(G1054_196_gat), .B(G1048_62_gat), .Y(G1063_242_gat) );
AND2XL U_g194 (.A(G1054_196_gat), .B(G200_25_gat), .Y(G1060_243_gat) );
AND2XL U_g195 (.A(G1022_206_gat), .B(G116_13_gat), .Y(G1025_244_gat) );
BUFX20 U_g196 (.A(G3040_152_gat), .Y(G3044_245_gat) );
AND2XL U_g197 (.A(G905_155_gat), .B(G540_65_gat), .Y(G630_246_gat) );
AND2XL U_g198 (.A(G905_155_gat), .B(G540_65_gat), .Y(G634_247_gat) );
AND2XL U_g199 (.A(G3101_160_gat), .B(G3098_153_gat), .Y(G646_248_gat) );
BUFX20 U_g200 (.A(G3098_153_gat), .Y(G3102_249_gat) );
AND2XL U_g201 (.A(G3109_159_gat), .B(G3106_154_gat), .Y(G912_250_gat) );
BUFX20 U_g202 (.A(G3106_154_gat), .Y(G3110_251_gat) );
AND2XL U_g203 (.A(G1001_203_gat), .B(G906_156_gat), .Y(G1004_252_gat) );
AND2XL U_g204 (.A(G1015_205_gat), .B(G851_68_gat), .Y(G1018_253_gat) );
BUFX20 U_g205 (.A(G3037_157_gat), .Y(G3043_254_gat) );
BUFX20 U_g206 (.A(G3030_161_gat), .Y(G3034_255_gat) );
AND2XL U_g207 (.A(G626_158_gat), .B(G87_10_gat), .Y(G654_256_gat) );
AND2XL U_g208 (.A(G626_158_gat), .B(G87_10_gat), .Y(G354_257_gat) );
BUFX20 U_g209 (.A(G3027_162_gat), .Y(G3033_258_gat) );
AND2XL U_g210 (.A(G994_202_gat), .B(G77_9_gat), .Y(G997_259_gat) );
AND2XL U_g211 (.A(G625_167_gat), .B(G479_82_gat), .Y(G352_260_gat) );
BUFX20 U_g212 (.A(G3020_163_gat), .Y(G3024_261_gat) );
AND2XL U_g213 (.A(G3085_172_gat), .B(G3082_165_gat), .Y(G642_262_gat) );
BUFX20 U_g214 (.A(G3082_165_gat), .Y(G3086_263_gat) );
AND2XL U_g215 (.A(G3093_171_gat), .B(G3090_166_gat), .Y(G903_264_gat) );
BUFX20 U_g216 (.A(G3090_166_gat), .Y(G3094_265_gat) );
AND2XL U_g217 (.A(G973_199_gat), .B(G897_168_gat), .Y(G976_266_gat) );
AND2XL U_g218 (.A(G987_201_gat), .B(G836_85_gat), .Y(G990_267_gat) );
BUFX20 U_g219 (.A(G3017_169_gat), .Y(G3023_268_gat) );
AND2XL U_g220 (.A(G636_175_gat), .B(G460_89_gat), .Y(G644_269_gat) );
AND2XL U_g221 (.A(G3013_174_gat), .B(G3010_173_gat), .Y(G3015_270_gat) );
BUFX20 U_g222 (.A(G3010_173_gat), .Y(G3014_271_gat) );
BUFX20 U_g223 (.A(G636_175_gat), .Y(G639_272_gat) );
AND2XL U_g224 (.A(G621_170_gat), .B(G432_99_gat), .Y(G650_273_gat) );
BUFX20 U_g225 (.A(G657_177_gat), .Y(G660_274_gat) );
BUFX20 U_g226 (.A(G675_178_gat), .Y(G678_275_gat) );
BUFX20 U_g227 (.A(G816_179_gat), .Y(G2128_276_gat) );
BUFX20 U_g228 (.A(G816_179_gat), .Y(G2181_277_gat) );
BUFX20 U_g229 (.A(G816_179_gat), .Y(G2233_278_gat) );
BUFX20 U_g230 (.A(G823_180_gat), .Y(G2076_279_gat) );
BUFX20 U_g231 (.A(G807_181_gat), .Y(G1870_280_gat) );
BUFX20 U_g232 (.A(G807_181_gat), .Y(G1920_281_gat) );
BUFX20 U_g233 (.A(G807_181_gat), .Y(G1971_282_gat) );
BUFX20 U_g234 (.A(G807_181_gat), .Y(G2021_283_gat) );
AND2XL U_g235 (.A(G794_182_gat), .B(G784_191_gat), .Y(G1527_284_gat) );
AND2XL U_g236 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1718_285_gat) );
AND2XL U_g237 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1725_286_gat) );
AND2XL U_g238 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1732_287_gat) );
AND2XL U_g239 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1739_288_gat) );
AND2XL U_g240 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1746_289_gat) );
AND2XL U_g241 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1753_290_gat) );
AND2XL U_g242 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1760_291_gat) );
AND2XL U_g243 (.A(G1699_105_gat), .B(G1681_192_gat), .Y(G1767_292_gat) );
AND2XL U_g244 (.A(G780_106_gat), .B(G860_208_gat), .Y(G806_293_gat) );
BUFX20 U_g245 (.A(G1681_192_gat), .Y(G1716_294_gat) );
BUFX20 U_g246 (.A(G1681_192_gat), .Y(G1723_295_gat) );
BUFX20 U_g247 (.A(G1681_192_gat), .Y(G1730_296_gat) );
BUFX20 U_g248 (.A(G1681_192_gat), .Y(G1737_297_gat) );
BUFX20 U_g249 (.A(G1681_192_gat), .Y(G1744_298_gat) );
BUFX20 U_g250 (.A(G1681_192_gat), .Y(G1751_299_gat) );
BUFX20 U_g251 (.A(G1681_192_gat), .Y(G1758_300_gat) );
BUFX20 U_g252 (.A(G1681_192_gat), .Y(G1765_301_gat) );
AND2XL U_g253 (.A(G794_182_gat), .B(G776_107_gat), .Y(G1530_302_gat) );
AND2XL U_g254 (.A(G776_107_gat), .B(G860_208_gat), .Y(G804_303_gat) );
BUFX20 U_g255 (.A(G1512_193_gat), .Y(G1581_304_gat) );
BUFX20 U_g256 (.A(G1512_193_gat), .Y(G1585_305_gat) );
BUFX20 U_g257 (.A(G1512_193_gat), .Y(G1589_306_gat) );
BUFX20 U_g258 (.A(G1512_193_gat), .Y(G1593_307_gat) );
BUFX20 U_g259 (.A(G1512_193_gat), .Y(G1597_308_gat) );
BUFX20 U_g260 (.A(G1512_193_gat), .Y(G1601_309_gat) );
BUFX20 U_g261 (.A(G1512_193_gat), .Y(G1605_310_gat) );
AND2XL U_g262 (.A(G1057_197_gat), .B(G1050_113_gat), .Y(G1069_311_gat) );
AND2XL U_g263 (.A(G1057_197_gat), .B(G1049_114_gat), .Y(G1066_312_gat) );
BUFX20 U_g264 (.A(G759_198_gat), .Y(G974_313_gat) );
BUFX20 U_g265 (.A(G759_198_gat), .Y(G981_314_gat) );
BUFX20 U_g266 (.A(G759_198_gat), .Y(G988_315_gat) );
BUFX20 U_g267 (.A(G759_198_gat), .Y(G995_316_gat) );
BUFX20 U_g268 (.A(G759_198_gat), .Y(G1002_317_gat) );
BUFX20 U_g269 (.A(G759_198_gat), .Y(G1009_318_gat) );
BUFX20 U_g270 (.A(G759_198_gat), .Y(G1016_319_gat) );
BUFX20 U_g271 (.A(G759_198_gat), .Y(G1023_320_gat) );
AND2XL U_g272 (.A(G759_198_gat), .B(G741_116_gat), .Y(G975_321_gat) );
AND2XL U_g273 (.A(G759_198_gat), .B(G741_116_gat), .Y(G982_322_gat) );
AND2XL U_g274 (.A(G759_198_gat), .B(G741_116_gat), .Y(G989_323_gat) );
AND2XL U_g275 (.A(G759_198_gat), .B(G741_116_gat), .Y(G996_324_gat) );
AND2XL U_g276 (.A(G759_198_gat), .B(G741_116_gat), .Y(G1003_325_gat) );
AND2XL U_g277 (.A(G759_198_gat), .B(G741_116_gat), .Y(G1010_326_gat) );
AND2XL U_g278 (.A(G759_198_gat), .B(G741_116_gat), .Y(G1017_327_gat) );
AND2XL U_g279 (.A(G759_198_gat), .B(G741_116_gat), .Y(G1024_328_gat) );
AND3XL U_g280 (.A(G784_191_gat), .B(G732_117_gat), .C(G724_119_gat), .Y(G1563_329_gat) );
AND3XL U_g281 (.A(G736_118_gat), .B(G721_211_gat), .C(G707_127_gat), .Y(G855_330_gat) );
BUFX20 U_g282 (.A(G861_209_gat), .Y(G915_331_gat) );
AND4XL U_g283 (.A(G794_182_gat), .B(G736_118_gat), .C(G724_119_gat), .D(G707_127_gat), .Y(G867_332_gat) );
BUFX20 U_g284 (.A(G864_210_gat), .Y(G941_333_gat) );
AND2XL U_g285 (.A(G784_191_gat), .B(G724_119_gat), .Y(G1572_334_gat) );
BUFX20 U_g286 (.A(G1834_215_gat), .Y(G1851_335_gat) );
BUFX20 U_g287 (.A(G1834_215_gat), .Y(G1901_336_gat) );
BUFX20 U_g288 (.A(G1834_215_gat), .Y(G1952_337_gat) );
BUFX20 U_g289 (.A(G1834_215_gat), .Y(G2002_338_gat) );
BUFX20 U_g290 (.A(G1834_215_gat), .Y(G2057_339_gat) );
BUFX20 U_g291 (.A(G1834_215_gat), .Y(G2109_340_gat) );
BUFX20 U_g292 (.A(G1834_215_gat), .Y(G2162_341_gat) );
BUFX20 U_g293 (.A(G1834_215_gat), .Y(G2214_342_gat) );
AND3XL U_g294 (.A(G1808_195_gat), .B(G13_1_gat), .C(G1_0_gat), .Y(G1809_343_gat) );
AND3XL U_g295 (.A(G1790_194_gat), .B(G13_1_gat), .C(G1_0_gat), .Y(G1791_344_gat) );
AND2XL U_g296 (.A(G1772_212_ngat), .B(G1_0_ngat), .Y(G1773_345_gat) );
AND2XL U_g297 (.A(G896_176_gat), .B(G890_125_gat), .Y(G956_346_gat) );
BUFX20 U_g298 (.A(G893_216_gat), .Y(G927_347_gat) );
AND3XL U_g299 (.A(G1541_151_gat), .B(G721_211_gat), .C(G707_127_gat), .Y(G1542_348_gat) );
AND2XL U_g300 (.A(G2897_49_gat), .B(G2877_217_gat), .Y(G2903_349_gat) );
AND2XL U_g301 (.A(G2897_49_gat), .B(G2877_217_gat), .Y(G2900_350_gat) );
AND2XL U_g302 (.A(G1765_301_gat), .B(G303_40_gat), .Y(G1768_351_gat) );
AND2XL U_g303 (.A(G1758_300_gat), .B(G294_39_gat), .Y(G1761_352_gat) );
AND2XL U_g304 (.A(G1751_299_gat), .B(G283_38_gat), .Y(G1754_353_gat) );
AND2XL U_g305 (.A(G1023_320_gat), .B(G283_38_gat), .Y(G1026_354_gat) );
AND2XL U_g306 (.A(G2966_220_gat), .B(G2965_218_gat), .Y(G2986_355_gat) );
AND2XL U_g307 (.A(G554_219_gat), .B(G553_227_gat), .Y(G586_356_gat) );
AND2XL U_g308 (.A(G1767_292_gat), .B(G264_35_gat), .Y(G1770_357_gat) );
AND2XL U_g309 (.A(G1760_291_gat), .B(G257_34_gat), .Y(G1763_358_gat) );
AND2XL U_g310 (.A(G2956_224_gat), .B(G2955_222_gat), .Y(G2983_359_gat) );
AND2XL U_g311 (.A(G1753_290_gat), .B(G250_33_gat), .Y(G1756_360_gat) );
AND2XL U_g312 (.A(G915_331_gat), .B(G588_137_gat), .Y(G920_361_gat) );
AND2XL U_g313 (.A(G1746_289_gat), .B(G244_32_gat), .Y(G1749_362_gat) );
AND2XL U_g314 (.A(G561_229_gat), .B(G560_226_gat), .Y(G562_363_gat) );
AND2XL U_g315 (.A(G1739_288_gat), .B(G238_31_gat), .Y(G1742_364_gat) );
AND2XL U_g316 (.A(G1732_287_gat), .B(G232_30_gat), .Y(G1735_365_gat) );
AND2XL U_g317 (.A(G556_233_gat), .B(G555_231_gat), .Y(G557_366_gat) );
AND2XL U_g318 (.A(G1725_286_gat), .B(G226_29_gat), .Y(G1728_367_gat) );
AND2XL U_g319 (.A(G1718_285_gat), .B(G223_28_gat), .Y(G1721_368_gat) );
BUFX20 U_g320 (.A(G2293_238_gat), .Y(G2485_369_gat) );
AND2XL U_g321 (.A(G1069_311_gat), .B(G1038_148_gat), .Y(G1096_370_gat) );
AND2XL U_g322 (.A(G1066_312_gat), .B(G1038_148_gat), .Y(G1108_371_gat) );
AND2XL U_g323 (.A(G1063_242_gat), .B(G1038_148_gat), .Y(G1144_372_gat) );
AND2XL U_g324 (.A(G1060_243_gat), .B(G1038_148_gat), .Y(G1156_373_gat) );
AND2XL U_g325 (.A(G1069_311_gat), .B(G1043_149_gat), .Y(G1072_374_gat) );
AND2XL U_g326 (.A(G1066_312_gat), .B(G1043_149_gat), .Y(G1084_375_gat) );
AND2XL U_g327 (.A(G1063_242_gat), .B(G1043_149_gat), .Y(G1120_376_gat) );
AND2XL U_g328 (.A(G1060_243_gat), .B(G1043_149_gat), .Y(G1132_377_gat) );
AND2XL U_g329 (.A(G982_322_gat), .B(G159_21_gat), .Y(G985_378_gat) );
AND2XL U_g330 (.A(G975_321_gat), .B(G150_20_gat), .Y(G978_379_gat) );
AND2XL U_g331 (.A(G1773_345_ngat), .B(G116_13_ngat), .Y(G2219_380_gat) );
AND2XL U_g332 (.A(G1744_298_gat), .B(G116_13_gat), .Y(G1747_381_gat) );
AND2XL U_g333 (.A(G1016_319_gat), .B(G116_13_gat), .Y(G1019_382_gat) );
AND2XL U_g334 (.A(G3043_254_gat), .B(G3040_152_gat), .Y(G3045_383_gat) );
AND2XL U_g335 (.A(G1773_345_ngat), .B(G107_12_ngat), .Y(G2167_384_gat) );
AND2XL U_g336 (.A(G1737_297_gat), .B(G107_12_gat), .Y(G1740_385_gat) );
AND2XL U_g337 (.A(G1009_318_gat), .B(G107_12_gat), .Y(G1012_386_gat) );
AND2XL U_g338 (.A(G3044_245_gat), .B(G3037_157_gat), .Y(G3046_387_gat) );
AND2XL U_g339 (.A(G1773_345_ngat), .B(G97_11_ngat), .Y(G2114_388_gat) );
AND2XL U_g340 (.A(G1730_296_gat), .B(G97_11_gat), .Y(G1733_389_gat) );
AND2XL U_g341 (.A(G3110_251_gat), .B(G3103_71_gat), .Y(G913_390_gat) );
AND2XL U_g342 (.A(G3102_249_gat), .B(G3095_72_gat), .Y(G647_391_gat) );
AND2XL U_g343 (.A(G1002_317_gat), .B(G845_74_gat), .Y(G1005_392_gat) );
AND2XL U_g344 (.A(G1024_328_gat), .B(G845_74_gat), .Y(G1027_393_gat) );
AND2XL U_g345 (.A(G3033_258_gat), .B(G3030_161_gat), .Y(G3035_394_gat) );
AND2XL U_g346 (.A(G1773_345_ngat), .B(G87_10_ngat), .Y(G2062_395_gat) );
AND2XL U_g347 (.A(G1723_295_gat), .B(G87_10_gat), .Y(G1726_396_gat) );
AND2XL U_g348 (.A(G995_316_gat), .B(G839_78_gat), .Y(G998_397_gat) );
AND2XL U_g349 (.A(G1017_327_gat), .B(G839_78_gat), .Y(G1020_398_gat) );
BUFX20 U_g350 (.A(G354_257_gat), .Y(G355_399_gat) );
AND2XL U_g351 (.A(G3034_255_gat), .B(G3027_162_gat), .Y(G3036_400_gat) );
AND2XL U_g352 (.A(G1773_345_ngat), .B(G77_9_ngat), .Y(G2007_401_gat) );
AND2XL U_g353 (.A(G1716_294_gat), .B(G77_9_gat), .Y(G1719_402_gat) );
AND2XL U_g354 (.A(G1010_326_gat), .B(G77_9_gat), .Y(G1013_403_gat) );
AND2XL U_g355 (.A(G988_315_gat), .B(G77_9_gat), .Y(G991_404_gat) );
BUFX20 U_g356 (.A(G352_260_gat), .Y(G353_405_gat) );
AND2XL U_g357 (.A(G3023_268_gat), .B(G3020_163_gat), .Y(G3025_406_gat) );
AND2XL U_g358 (.A(G1773_345_ngat), .B(G68_8_ngat), .Y(G1957_407_gat) );
AND2XL U_g359 (.A(G981_314_gat), .B(G833_86_gat), .Y(G984_408_gat) );
AND2XL U_g360 (.A(G1003_325_gat), .B(G833_86_gat), .Y(G1006_409_gat) );
AND2XL U_g361 (.A(G3024_261_gat), .B(G3017_169_gat), .Y(G3026_410_gat) );
AND2XL U_g362 (.A(G1773_345_ngat), .B(G58_7_ngat), .Y(G1906_411_gat) );
AND2XL U_g363 (.A(G3094_265_gat), .B(G3087_90_gat), .Y(G904_412_gat) );
AND2XL U_g364 (.A(G3086_263_gat), .B(G3079_91_gat), .Y(G643_413_gat) );
AND2XL U_g365 (.A(G974_313_gat), .B(G828_93_gat), .Y(G977_414_gat) );
AND2XL U_g366 (.A(G996_324_gat), .B(G828_93_gat), .Y(G999_415_gat) );
AND4XL U_g367 (.A(G58_7_gat), .B(G442_98_gat), .C(G635_164_gat), .D(G630_246_gat), .Y(G655_416_gat) );
AND2XL U_g368 (.A(G1773_345_ngat), .B(G50_6_ngat), .Y(G1856_417_gat) );
AND2XL U_g369 (.A(G989_323_gat), .B(G50_6_gat), .Y(G992_418_gat) );
AND2XL U_g370 (.A(G3014_271_gat), .B(G3007_97_gat), .Y(G3016_419_gat) );
AND2XL U_g371 (.A(G675_178_gat), .B(G650_273_gat), .Y(G680_420_gat) );
BUFX20 U_g372 (.A(G1527_284_gat), .Y(G1533_421_gat) );
AND2XL U_g373 (.A(G1530_302_gat), .B(G1527_284_gat), .Y(G1535_422_gat) );
AND2XL U_g374 (.A(G806_293_gat), .B(G804_303_gat), .Y(G613_423_gat) );
BUFX20 U_g375 (.A(G806_293_gat), .Y(G616_424_gat) );
AND2XL U_g376 (.A(G806_293_gat), .B(G804_303_gat), .Y(G668_425_gat) );
BUFX20 U_g377 (.A(G806_293_gat), .Y(G671_426_gat) );
BUFX20 U_g378 (.A(G806_293_gat), .Y(G685_427_gat) );
AND2XL U_g379 (.A(G806_293_gat), .B(G804_303_gat), .Y(G688_428_gat) );
BUFX20 U_g380 (.A(G806_293_gat), .Y(G696_429_gat) );
AND2XL U_g381 (.A(G806_293_gat), .B(G804_303_gat), .Y(G699_430_gat) );
BUFX20 U_g382 (.A(G1530_302_gat), .Y(G1534_431_gat) );
BUFX20 U_g383 (.A(G804_303_gat), .Y(G610_432_gat) );
BUFX20 U_g384 (.A(G804_303_gat), .Y(G665_433_gat) );
BUFX20 U_g385 (.A(G804_303_gat), .Y(G683_434_gat) );
BUFX20 U_g386 (.A(G804_303_gat), .Y(G694_435_gat) );
BUFX20 U_g387 (.A(G1563_329_gat), .Y(G1646_436_gat) );
BUFX20 U_g388 (.A(G1563_329_gat), .Y(G1655_437_gat) );
BUFX20 U_g389 (.A(G1563_329_gat), .Y(G1664_438_gat) );
BUFX20 U_g390 (.A(G1563_329_gat), .Y(G1673_439_gat) );
BUFX20 U_g391 (.A(G855_330_gat), .Y(G914_440_gat) );
BUFX20 U_g392 (.A(G855_330_gat), .Y(G942_441_gat) );
AND2XL U_g393 (.A(G861_209_gat), .B(G855_330_gat), .Y(G916_442_gat) );
BUFX20 U_g394 (.A(G867_332_gat), .Y(G870_443_gat) );
BUFX20 U_g395 (.A(G867_332_gat), .Y(G887_444_gat) );
AND2XL U_g396 (.A(G855_330_gat), .B(G864_210_gat), .Y(G943_445_gat) );
BUFX20 U_g397 (.A(G1572_334_gat), .Y(G1610_446_gat) );
BUFX20 U_g398 (.A(G1572_334_gat), .Y(G1619_447_gat) );
BUFX20 U_g399 (.A(G1572_334_gat), .Y(G1628_448_gat) );
BUFX20 U_g400 (.A(G1572_334_gat), .Y(G1637_449_gat) );
AND2XL U_g401 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G1852_450_gat) );
AND2XL U_g402 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G1902_451_gat) );
AND2XL U_g403 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G1953_452_gat) );
AND2XL U_g404 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G2003_453_gat) );
AND2XL U_g405 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G2058_454_gat) );
AND2XL U_g406 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G2110_455_gat) );
AND2XL U_g407 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G2163_456_gat) );
AND2XL U_g408 (.A(G1773_345_gat), .B(G1834_215_gat), .Y(G2215_457_gat) );
BUFX20 U_g409 (.A(G1809_343_gat), .Y(G1812_458_gat) );
BUFX20 U_g410 (.A(G1809_343_gat), .Y(G1817_459_gat) );
BUFX20 U_g411 (.A(G1791_344_gat), .Y(G1794_460_gat) );
BUFX20 U_g412 (.A(G1791_344_gat), .Y(G1799_461_gat) );
BUFX20 U_g413 (.A(G956_346_gat), .Y(G2678_462_gat) );
BUFX20 U_g414 (.A(G956_346_gat), .Y(G2697_463_gat) );
BUFX20 U_g415 (.A(G956_346_gat), .Y(G2716_464_gat) );
BUFX20 U_g416 (.A(G956_346_gat), .Y(G2733_465_gat) );
BUFX20 U_g417 (.A(G956_346_gat), .Y(G2751_466_gat) );
BUFX20 U_g418 (.A(G956_346_gat), .Y(G2768_467_gat) );
BUFX20 U_g419 (.A(G956_346_gat), .Y(G2785_468_gat) );
BUFX20 U_g420 (.A(G956_346_gat), .Y(G2802_469_gat) );
BUFX20 U_g421 (.A(G1542_348_gat), .Y(G1545_470_gat) );
BUFX20 U_g422 (.A(G1542_348_gat), .Y(G1554_471_gat) );
AND3XL U_g423 (.A(G816_179_gat), .B(G274_37_gat), .C(G1799_461_gat), .Y(G2235_472_gat) );
AND3XL U_g424 (.A(G816_179_gat), .B(G274_37_gat), .C(G1799_461_gat), .Y(G2183_473_gat) );
AND3XL U_g425 (.A(G816_179_gat), .B(G274_37_gat), .C(G1799_461_gat), .Y(G2130_474_gat) );
AND3XL U_g426 (.A(G823_180_gat), .B(G274_37_gat), .C(G1799_461_gat), .Y(G2078_475_gat) );
AND3XL U_g427 (.A(G807_181_gat), .B(G274_37_gat), .C(G1817_459_gat), .Y(G2023_476_gat) );
AND3XL U_g428 (.A(G807_181_gat), .B(G274_37_gat), .C(G1817_459_gat), .Y(G1973_477_gat) );
AND3XL U_g429 (.A(G807_181_gat), .B(G274_37_gat), .C(G1817_459_gat), .Y(G1922_478_gat) );
AND3XL U_g430 (.A(G807_181_gat), .B(G274_37_gat), .C(G1817_459_gat), .Y(G1872_479_gat) );
AND3XL U_g431 (.A(G2233_278_gat), .B(G270_36_gat), .C(G1799_461_gat), .Y(G2234_480_gat) );
BUFX20 U_g432 (.A(G2986_355_gat), .Y(G2990_481_gat) );
AND2XL U_g433 (.A(G916_442_gat), .B(G586_356_gat), .Y(G923_482_gat) );
AND3XL U_g434 (.A(G2181_277_gat), .B(G264_35_gat), .C(G1799_461_gat), .Y(G2182_483_gat) );
AND3XL U_g435 (.A(G2128_276_gat), .B(G257_34_gat), .C(G1799_461_gat), .Y(G2129_484_gat) );
AND3XL U_g436 (.A(G1770_357_ngat), .B(G1769_221_ngat), .C(G1768_351_ngat), .Y(G1771_485_gat) );
BUFX20 U_g437 (.A(G2983_359_gat), .Y(G2989_486_gat) );
AND3XL U_g438 (.A(G2076_279_gat), .B(G250_33_gat), .C(G1799_461_gat), .Y(G2077_487_gat) );
AND3XL U_g439 (.A(G1763_358_ngat), .B(G1762_223_ngat), .C(G1761_352_ngat), .Y(G1764_488_gat) );
AND3XL U_g440 (.A(G2021_283_gat), .B(G244_32_gat), .C(G1817_459_gat), .Y(G2022_489_gat) );
AND3XL U_g441 (.A(G1756_360_ngat), .B(G1755_225_ngat), .C(G1754_353_ngat), .Y(G1757_490_gat) );
BUFX20 U_g442 (.A(G562_363_gat), .Y(G2970_491_gat) );
BUFX20 U_g443 (.A(G562_363_gat), .Y(G2978_492_gat) );
AND3XL U_g444 (.A(G1971_282_gat), .B(G238_31_gat), .C(G1817_459_gat), .Y(G1972_493_gat) );
AND3XL U_g445 (.A(G1749_362_ngat), .B(G1748_228_ngat), .C(G1747_381_ngat), .Y(G1750_494_gat) );
AND3XL U_g446 (.A(G1920_281_gat), .B(G232_30_gat), .C(G1817_459_gat), .Y(G1921_495_gat) );
AND3XL U_g447 (.A(G1742_364_ngat), .B(G1741_230_ngat), .C(G1740_385_ngat), .Y(G1743_496_gat) );
BUFX20 U_g448 (.A(G557_366_gat), .Y(G2967_497_gat) );
BUFX20 U_g449 (.A(G557_366_gat), .Y(G2975_498_gat) );
AND3XL U_g450 (.A(G1870_280_gat), .B(G226_29_gat), .C(G1817_459_gat), .Y(G1871_499_gat) );
AND3XL U_g451 (.A(G1735_365_ngat), .B(G1734_232_ngat), .C(G1733_389_ngat), .Y(G1736_500_gat) );
AND3XL U_g452 (.A(G1728_367_ngat), .B(G1727_234_ngat), .C(G1726_396_ngat), .Y(G1729_501_gat) );
AND3XL U_g453 (.A(G1721_368_ngat), .B(G1720_235_ngat), .C(G1719_402_ngat), .Y(G1722_502_gat) );
BUFX20 U_g454 (.A(G2485_369_gat), .Y(G2488_503_gat) );
BUFX20 U_g455 (.A(G1096_370_gat), .Y(G1099_504_gat) );
BUFX20 U_g456 (.A(G1096_370_gat), .Y(G1186_505_gat) );
BUFX20 U_g457 (.A(G1108_371_gat), .Y(G1111_506_gat) );
BUFX20 U_g458 (.A(G1108_371_gat), .Y(G1195_507_gat) );
BUFX20 U_g459 (.A(G1144_372_gat), .Y(G1147_508_gat) );
BUFX20 U_g460 (.A(G1144_372_gat), .Y(G1222_509_gat) );
BUFX20 U_g461 (.A(G1156_373_gat), .Y(G1159_510_gat) );
BUFX20 U_g462 (.A(G1156_373_gat), .Y(G1231_511_gat) );
BUFX20 U_g463 (.A(G1072_374_gat), .Y(G1075_512_gat) );
BUFX20 U_g464 (.A(G1072_374_gat), .Y(G1168_513_gat) );
BUFX20 U_g465 (.A(G1084_375_gat), .Y(G1087_514_gat) );
BUFX20 U_g466 (.A(G1084_375_gat), .Y(G1177_515_gat) );
BUFX20 U_g467 (.A(G1120_376_gat), .Y(G1123_516_gat) );
BUFX20 U_g468 (.A(G1120_376_gat), .Y(G1204_517_gat) );
BUFX20 U_g469 (.A(G1132_377_gat), .Y(G1135_518_gat) );
BUFX20 U_g470 (.A(G1132_377_gat), .Y(G1213_519_gat) );
AND3XL U_g471 (.A(G2215_457_gat), .B(G2052_213_gat), .C(G116_13_gat), .Y(G2222_520_gat) );
AND3XL U_g472 (.A(G1027_393_ngat), .B(G1026_354_ngat), .C(G1025_244_ngat), .Y(G1028_521_gat) );
AND2XL U_g473 (.A(G3046_387_gat), .B(G3045_383_gat), .Y(G3058_522_gat) );
AND2XL U_g474 (.A(G696_429_gat), .B(G634_247_gat), .Y(G701_523_gat) );
AND2XL U_g475 (.A(G688_428_gat), .B(G540_65_gat), .Y(G691_524_gat) );
AND3XL U_g476 (.A(G2163_456_gat), .B(G2052_213_gat), .C(G107_12_gat), .Y(G2170_525_gat) );
AND2XL U_g477 (.A(G647_391_gat), .B(G646_248_gat), .Y(G648_526_gat) );
AND2XL U_g478 (.A(G913_390_gat), .B(G912_250_gat), .Y(G910_527_gat) );
AND3XL U_g479 (.A(G1006_409_ngat), .B(G1005_392_ngat), .C(G1004_252_ngat), .Y(G1007_528_gat) );
AND3XL U_g480 (.A(G1020_398_ngat), .B(G1019_382_ngat), .C(G1018_253_ngat), .Y(G1021_529_gat) );
AND2XL U_g481 (.A(G699_430_gat), .B(G526_69_gat), .Y(G702_530_gat) );
AND3XL U_g482 (.A(G2110_455_gat), .B(G2052_213_gat), .C(G97_11_gat), .Y(G2117_531_gat) );
AND2XL U_g483 (.A(G3036_400_gat), .B(G3035_394_gat), .Y(G3055_532_gat) );
AND2XL U_g484 (.A(G668_425_gat), .B(G513_75_gat), .Y(G672_533_gat) );
AND3XL U_g485 (.A(G2058_454_gat), .B(G2052_213_gat), .C(G87_10_gat), .Y(G2065_534_gat) );
AND2XL U_g486 (.A(G685_427_gat), .B(G654_256_gat), .Y(G690_535_gat) );
AND2XL U_g487 (.A(G613_423_gat), .B(G501_79_gat), .Y(G617_536_gat) );
AND3XL U_g488 (.A(G2003_453_gat), .B(G1829_214_gat), .C(G77_9_gat), .Y(G2010_537_gat) );
AND3XL U_g489 (.A(G999_415_ngat), .B(G998_397_ngat), .C(G997_259_ngat), .Y(G1000_538_gat) );
AND2XL U_g490 (.A(G3026_410_gat), .B(G3025_406_gat), .Y(G3050_539_gat) );
AND3XL U_g491 (.A(G1953_452_gat), .B(G1829_214_gat), .C(G68_8_gat), .Y(G1960_540_gat) );
AND2XL U_g492 (.A(G643_413_gat), .B(G642_262_gat), .Y(G640_541_gat) );
AND2XL U_g493 (.A(G904_412_gat), .B(G903_264_gat), .Y(G901_542_gat) );
AND3XL U_g494 (.A(G978_379_ngat), .B(G977_414_ngat), .C(G976_266_ngat), .Y(G979_543_gat) );
AND3XL U_g495 (.A(G992_418_ngat), .B(G991_404_ngat), .C(G990_267_ngat), .Y(G993_544_gat) );
AND3XL U_g496 (.A(G1902_451_gat), .B(G1829_214_gat), .C(G58_7_gat), .Y(G1909_545_gat) );
AND2XL U_g497 (.A(G3016_419_gat), .B(G3015_270_gat), .Y(G3047_546_gat) );
AND3XL U_g498 (.A(G1852_450_gat), .B(G1829_214_gat), .C(G50_6_gat), .Y(G1859_547_gat) );
AND2XL U_g499 (.A(G1535_422_gat), .B(G442_98_gat), .Y(G1538_548_gat) );
AND2XL U_g500 (.A(G914_440_gat), .B(G650_273_gat), .Y(G917_549_gat) );
AND2XL U_g501 (.A(G657_177_gat), .B(G655_416_gat), .Y(G662_550_gat) );
AND2XL U_g502 (.A(G1563_329_gat), .B(G1554_471_gat), .Y(G1647_551_gat) );
AND2XL U_g503 (.A(G1563_329_gat), .B(G1554_471_gat), .Y(G1656_552_gat) );
AND2XL U_g504 (.A(G1563_329_gat), .B(G1554_471_gat), .Y(G1665_553_gat) );
AND2XL U_g505 (.A(G1563_329_gat), .B(G1554_471_gat), .Y(G1674_554_gat) );
BUFX20 U_g506 (.A(G870_443_gat), .Y(G2679_555_gat) );
BUFX20 U_g507 (.A(G870_443_gat), .Y(G2698_556_gat) );
BUFX20 U_g508 (.A(G870_443_gat), .Y(G2717_557_gat) );
BUFX20 U_g509 (.A(G870_443_gat), .Y(G2734_558_gat) );
BUFX20 U_g510 (.A(G870_443_gat), .Y(G2752_559_gat) );
BUFX20 U_g511 (.A(G870_443_gat), .Y(G2769_560_gat) );
BUFX20 U_g512 (.A(G870_443_gat), .Y(G2786_561_gat) );
BUFX20 U_g513 (.A(G870_443_gat), .Y(G2803_562_gat) );
BUFX20 U_g514 (.A(G887_444_gat), .Y(G926_563_gat) );
AND2XL U_g515 (.A(G1572_334_gat), .B(G1545_470_gat), .Y(G1611_564_gat) );
AND2XL U_g516 (.A(G1572_334_gat), .B(G1545_470_gat), .Y(G1620_565_gat) );
AND2XL U_g517 (.A(G1572_334_gat), .B(G1545_470_gat), .Y(G1629_566_gat) );
AND2XL U_g518 (.A(G1572_334_gat), .B(G1545_470_gat), .Y(G1638_567_gat) );
AND2XL U_g519 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2680_568_gat) );
AND2XL U_g520 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2699_569_gat) );
AND2XL U_g521 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2718_570_gat) );
AND2XL U_g522 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2735_571_gat) );
AND2XL U_g523 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2753_572_gat) );
AND2XL U_g524 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2770_573_gat) );
AND2XL U_g525 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2787_574_gat) );
AND2XL U_g526 (.A(G870_443_gat), .B(G956_346_gat), .Y(G2804_575_gat) );
AND2XL U_g527 (.A(G893_216_gat), .B(G887_444_gat), .Y(G928_576_gat) );
BUFX20 U_g528 (.A(G1545_470_gat), .Y(G1609_577_gat) );
BUFX20 U_g529 (.A(G1545_470_gat), .Y(G1618_578_gat) );
BUFX20 U_g530 (.A(G1545_470_gat), .Y(G1627_579_gat) );
BUFX20 U_g531 (.A(G1545_470_gat), .Y(G1636_580_gat) );
BUFX20 U_g532 (.A(G1554_471_gat), .Y(G1645_581_gat) );
BUFX20 U_g533 (.A(G1554_471_gat), .Y(G1654_582_gat) );
BUFX20 U_g534 (.A(G1554_471_gat), .Y(G1663_583_gat) );
BUFX20 U_g535 (.A(G1554_471_gat), .Y(G1672_584_gat) );
AND2XL U_g536 (.A(G2989_486_gat), .B(G2986_355_gat), .Y(G574_585_gat) );
AND2XL U_g537 (.A(G2990_481_gat), .B(G2983_359_gat), .Y(G575_586_gat) );
AND3XL U_g538 (.A(G923_482_ngat), .B(G920_361_ngat), .C(G917_549_ngat), .Y(G359_587_gat) );
AND3XL U_g539 (.A(G923_482_ngat), .B(G920_361_ngat), .C(G917_549_ngat), .Y(G1029_588_gat) );
BUFX20 U_g540 (.A(G2970_491_gat), .Y(G2974_589_gat) );
BUFX20 U_g541 (.A(G2978_492_gat), .Y(G2982_590_gat) );
BUFX20 U_g542 (.A(G2967_497_gat), .Y(G2973_591_gat) );
BUFX20 U_g543 (.A(G2975_498_gat), .Y(G2981_592_gat) );
BUFX20 U_g544 (.A(G1099_504_gat), .Y(G1242_593_gat) );
BUFX20 U_g545 (.A(G1099_504_gat), .Y(G1259_594_gat) );
BUFX20 U_g546 (.A(G1099_504_gat), .Y(G1276_595_gat) );
BUFX20 U_g547 (.A(G1099_504_gat), .Y(G1293_596_gat) );
BUFX20 U_g548 (.A(G1099_504_gat), .Y(G1310_597_gat) );
BUFX20 U_g549 (.A(G1099_504_gat), .Y(G1327_598_gat) );
BUFX20 U_g550 (.A(G1099_504_gat), .Y(G1344_599_gat) );
BUFX20 U_g551 (.A(G1099_504_gat), .Y(G1361_600_gat) );
BUFX20 U_g552 (.A(G1186_505_gat), .Y(G1378_601_gat) );
BUFX20 U_g553 (.A(G1186_505_gat), .Y(G1395_602_gat) );
BUFX20 U_g554 (.A(G1186_505_gat), .Y(G1412_603_gat) );
BUFX20 U_g555 (.A(G1186_505_gat), .Y(G1429_604_gat) );
BUFX20 U_g556 (.A(G1186_505_gat), .Y(G1446_605_gat) );
BUFX20 U_g557 (.A(G1186_505_gat), .Y(G1463_606_gat) );
BUFX20 U_g558 (.A(G1186_505_gat), .Y(G1480_607_gat) );
BUFX20 U_g559 (.A(G1186_505_gat), .Y(G1497_608_gat) );
BUFX20 U_g560 (.A(G1111_506_gat), .Y(G1243_609_gat) );
BUFX20 U_g561 (.A(G1111_506_gat), .Y(G1260_610_gat) );
BUFX20 U_g562 (.A(G1111_506_gat), .Y(G1277_611_gat) );
BUFX20 U_g563 (.A(G1111_506_gat), .Y(G1294_612_gat) );
BUFX20 U_g564 (.A(G1111_506_gat), .Y(G1311_613_gat) );
BUFX20 U_g565 (.A(G1111_506_gat), .Y(G1328_614_gat) );
BUFX20 U_g566 (.A(G1111_506_gat), .Y(G1345_615_gat) );
BUFX20 U_g567 (.A(G1111_506_gat), .Y(G1362_616_gat) );
BUFX20 U_g568 (.A(G1195_507_gat), .Y(G1379_617_gat) );
BUFX20 U_g569 (.A(G1195_507_gat), .Y(G1396_618_gat) );
BUFX20 U_g570 (.A(G1195_507_gat), .Y(G1413_619_gat) );
BUFX20 U_g571 (.A(G1195_507_gat), .Y(G1430_620_gat) );
BUFX20 U_g572 (.A(G1195_507_gat), .Y(G1447_621_gat) );
BUFX20 U_g573 (.A(G1195_507_gat), .Y(G1464_622_gat) );
BUFX20 U_g574 (.A(G1195_507_gat), .Y(G1481_623_gat) );
BUFX20 U_g575 (.A(G1195_507_gat), .Y(G1498_624_gat) );
BUFX20 U_g576 (.A(G1147_508_gat), .Y(G1246_625_gat) );
BUFX20 U_g577 (.A(G1147_508_gat), .Y(G1263_626_gat) );
BUFX20 U_g578 (.A(G1147_508_gat), .Y(G1280_627_gat) );
BUFX20 U_g579 (.A(G1147_508_gat), .Y(G1297_628_gat) );
BUFX20 U_g580 (.A(G1147_508_gat), .Y(G1314_629_gat) );
BUFX20 U_g581 (.A(G1147_508_gat), .Y(G1331_630_gat) );
BUFX20 U_g582 (.A(G1147_508_gat), .Y(G1348_631_gat) );
BUFX20 U_g583 (.A(G1147_508_gat), .Y(G1365_632_gat) );
BUFX20 U_g584 (.A(G1222_509_gat), .Y(G1382_633_gat) );
BUFX20 U_g585 (.A(G1222_509_gat), .Y(G1399_634_gat) );
BUFX20 U_g586 (.A(G1222_509_gat), .Y(G1416_635_gat) );
BUFX20 U_g587 (.A(G1222_509_gat), .Y(G1433_636_gat) );
BUFX20 U_g588 (.A(G1222_509_gat), .Y(G1450_637_gat) );
BUFX20 U_g589 (.A(G1222_509_gat), .Y(G1467_638_gat) );
BUFX20 U_g590 (.A(G1222_509_gat), .Y(G1484_639_gat) );
BUFX20 U_g591 (.A(G1222_509_gat), .Y(G1501_640_gat) );
BUFX20 U_g592 (.A(G1159_510_gat), .Y(G1247_641_gat) );
BUFX20 U_g593 (.A(G1159_510_gat), .Y(G1264_642_gat) );
BUFX20 U_g594 (.A(G1159_510_gat), .Y(G1281_643_gat) );
BUFX20 U_g595 (.A(G1159_510_gat), .Y(G1298_644_gat) );
BUFX20 U_g596 (.A(G1159_510_gat), .Y(G1315_645_gat) );
BUFX20 U_g597 (.A(G1159_510_gat), .Y(G1332_646_gat) );
BUFX20 U_g598 (.A(G1159_510_gat), .Y(G1349_647_gat) );
BUFX20 U_g599 (.A(G1159_510_gat), .Y(G1366_648_gat) );
BUFX20 U_g600 (.A(G1231_511_gat), .Y(G1383_649_gat) );
BUFX20 U_g601 (.A(G1231_511_gat), .Y(G1400_650_gat) );
BUFX20 U_g602 (.A(G1231_511_gat), .Y(G1417_651_gat) );
BUFX20 U_g603 (.A(G1231_511_gat), .Y(G1434_652_gat) );
BUFX20 U_g604 (.A(G1231_511_gat), .Y(G1451_653_gat) );
BUFX20 U_g605 (.A(G1231_511_gat), .Y(G1468_654_gat) );
BUFX20 U_g606 (.A(G1231_511_gat), .Y(G1485_655_gat) );
BUFX20 U_g607 (.A(G1231_511_gat), .Y(G1502_656_gat) );
BUFX20 U_g608 (.A(G1075_512_gat), .Y(G1240_657_gat) );
BUFX20 U_g609 (.A(G1075_512_gat), .Y(G1257_658_gat) );
BUFX20 U_g610 (.A(G1075_512_gat), .Y(G1274_659_gat) );
BUFX20 U_g611 (.A(G1075_512_gat), .Y(G1291_660_gat) );
BUFX20 U_g612 (.A(G1075_512_gat), .Y(G1308_661_gat) );
BUFX20 U_g613 (.A(G1075_512_gat), .Y(G1325_662_gat) );
BUFX20 U_g614 (.A(G1075_512_gat), .Y(G1342_663_gat) );
BUFX20 U_g615 (.A(G1075_512_gat), .Y(G1359_664_gat) );
BUFX20 U_g616 (.A(G1168_513_gat), .Y(G1376_665_gat) );
BUFX20 U_g617 (.A(G1168_513_gat), .Y(G1393_666_gat) );
BUFX20 U_g618 (.A(G1168_513_gat), .Y(G1410_667_gat) );
BUFX20 U_g619 (.A(G1168_513_gat), .Y(G1427_668_gat) );
BUFX20 U_g620 (.A(G1168_513_gat), .Y(G1444_669_gat) );
BUFX20 U_g621 (.A(G1168_513_gat), .Y(G1461_670_gat) );
BUFX20 U_g622 (.A(G1168_513_gat), .Y(G1478_671_gat) );
BUFX20 U_g623 (.A(G1168_513_gat), .Y(G1495_672_gat) );
BUFX20 U_g624 (.A(G1087_514_gat), .Y(G1241_673_gat) );
BUFX20 U_g625 (.A(G1087_514_gat), .Y(G1258_674_gat) );
BUFX20 U_g626 (.A(G1087_514_gat), .Y(G1275_675_gat) );
BUFX20 U_g627 (.A(G1087_514_gat), .Y(G1292_676_gat) );
BUFX20 U_g628 (.A(G1087_514_gat), .Y(G1309_677_gat) );
BUFX20 U_g629 (.A(G1087_514_gat), .Y(G1326_678_gat) );
BUFX20 U_g630 (.A(G1087_514_gat), .Y(G1343_679_gat) );
BUFX20 U_g631 (.A(G1087_514_gat), .Y(G1360_680_gat) );
BUFX20 U_g632 (.A(G1177_515_gat), .Y(G1377_681_gat) );
BUFX20 U_g633 (.A(G1177_515_gat), .Y(G1394_682_gat) );
BUFX20 U_g634 (.A(G1177_515_gat), .Y(G1411_683_gat) );
BUFX20 U_g635 (.A(G1177_515_gat), .Y(G1428_684_gat) );
BUFX20 U_g636 (.A(G1177_515_gat), .Y(G1445_685_gat) );
BUFX20 U_g637 (.A(G1177_515_gat), .Y(G1462_686_gat) );
BUFX20 U_g638 (.A(G1177_515_gat), .Y(G1479_687_gat) );
BUFX20 U_g639 (.A(G1177_515_gat), .Y(G1496_688_gat) );
BUFX20 U_g640 (.A(G1123_516_gat), .Y(G1244_689_gat) );
BUFX20 U_g641 (.A(G1123_516_gat), .Y(G1261_690_gat) );
BUFX20 U_g642 (.A(G1123_516_gat), .Y(G1278_691_gat) );
BUFX20 U_g643 (.A(G1123_516_gat), .Y(G1295_692_gat) );
BUFX20 U_g644 (.A(G1123_516_gat), .Y(G1312_693_gat) );
BUFX20 U_g645 (.A(G1123_516_gat), .Y(G1329_694_gat) );
BUFX20 U_g646 (.A(G1123_516_gat), .Y(G1346_695_gat) );
BUFX20 U_g647 (.A(G1123_516_gat), .Y(G1363_696_gat) );
BUFX20 U_g648 (.A(G1204_517_gat), .Y(G1380_697_gat) );
BUFX20 U_g649 (.A(G1204_517_gat), .Y(G1397_698_gat) );
BUFX20 U_g650 (.A(G1204_517_gat), .Y(G1414_699_gat) );
BUFX20 U_g651 (.A(G1204_517_gat), .Y(G1431_700_gat) );
BUFX20 U_g652 (.A(G1204_517_gat), .Y(G1448_701_gat) );
BUFX20 U_g653 (.A(G1204_517_gat), .Y(G1465_702_gat) );
BUFX20 U_g654 (.A(G1204_517_gat), .Y(G1482_703_gat) );
BUFX20 U_g655 (.A(G1204_517_gat), .Y(G1499_704_gat) );
BUFX20 U_g656 (.A(G1135_518_gat), .Y(G1245_705_gat) );
BUFX20 U_g657 (.A(G1135_518_gat), .Y(G1262_706_gat) );
BUFX20 U_g658 (.A(G1135_518_gat), .Y(G1279_707_gat) );
BUFX20 U_g659 (.A(G1135_518_gat), .Y(G1296_708_gat) );
BUFX20 U_g660 (.A(G1135_518_gat), .Y(G1313_709_gat) );
BUFX20 U_g661 (.A(G1135_518_gat), .Y(G1330_710_gat) );
BUFX20 U_g662 (.A(G1135_518_gat), .Y(G1347_711_gat) );
BUFX20 U_g663 (.A(G1135_518_gat), .Y(G1364_712_gat) );
BUFX20 U_g664 (.A(G1213_519_gat), .Y(G1381_713_gat) );
BUFX20 U_g665 (.A(G1213_519_gat), .Y(G1398_714_gat) );
BUFX20 U_g666 (.A(G1213_519_gat), .Y(G1415_715_gat) );
BUFX20 U_g667 (.A(G1213_519_gat), .Y(G1432_716_gat) );
BUFX20 U_g668 (.A(G1213_519_gat), .Y(G1449_717_gat) );
BUFX20 U_g669 (.A(G1213_519_gat), .Y(G1466_718_gat) );
BUFX20 U_g670 (.A(G1213_519_gat), .Y(G1483_719_gat) );
BUFX20 U_g671 (.A(G1213_519_gat), .Y(G1500_720_gat) );
BUFX20 U_g672 (.A(G3058_522_gat), .Y(G3062_721_gat) );
AND2XL U_g673 (.A(G928_576_gat), .B(G630_246_gat), .Y(G938_722_gat) );
AND2XL U_g674 (.A(G648_526_gat), .B(G530_66_gat), .Y(G649_723_gat) );
BUFX20 U_g675 (.A(G910_527_gat), .Y(G911_724_gat) );
BUFX20 U_g676 (.A(G3055_532_gat), .Y(G3061_725_gat) );
BUFX20 U_g677 (.A(G3050_539_gat), .Y(G3054_726_gat) );
AND2XL U_g678 (.A(G1638_567_gat), .B(G479_82_gat), .Y(G1643_727_gat) );
AND3XL U_g679 (.A(G639_272_gat), .B(G476_83_gat), .C(G640_541_gat), .Y(G641_728_gat) );
BUFX20 U_g680 (.A(G901_542_gat), .Y(G902_729_gat) );
AND2XL U_g681 (.A(G1629_566_gat), .B(G463_88_gat), .Y(G1634_730_gat) );
BUFX20 U_g682 (.A(G3047_546_gat), .Y(G3053_731_gat) );
AND2XL U_g683 (.A(G1620_565_gat), .B(G456_94_gat), .Y(G1625_732_gat) );
AND2XL U_g684 (.A(G1611_564_gat), .B(G442_98_gat), .Y(G1616_733_gat) );
AND2XL U_g685 (.A(G926_563_gat), .B(G650_273_gat), .Y(G929_734_gat) );
AND2XL U_g686 (.A(G1851_335_gat), .B(G979_543_gat), .Y(G1853_735_gat) );
AND2XL U_g687 (.A(G1952_337_gat), .B(G993_544_gat), .Y(G1954_736_gat) );
AND2XL U_g688 (.A(G2002_338_gat), .B(G1000_538_gat), .Y(G2004_737_gat) );
AND2XL U_g689 (.A(G2057_339_gat), .B(G1007_528_gat), .Y(G2059_738_gat) );
AND2XL U_g690 (.A(G2162_341_gat), .B(G1021_529_gat), .Y(G2164_739_gat) );
AND2XL U_g691 (.A(G2214_342_gat), .B(G1028_521_gat), .Y(G2216_740_gat) );
AND2XL U_g692 (.A(G1722_502_gat), .B(G1812_458_gat), .Y(G1873_741_gat) );
AND2XL U_g693 (.A(G1729_501_gat), .B(G1812_458_gat), .Y(G1923_742_gat) );
AND2XL U_g694 (.A(G1736_500_gat), .B(G1812_458_gat), .Y(G1974_743_gat) );
AND2XL U_g695 (.A(G1743_496_gat), .B(G1812_458_gat), .Y(G2024_744_gat) );
AND2XL U_g696 (.A(G1750_494_gat), .B(G1794_460_gat), .Y(G2079_745_gat) );
AND2XL U_g697 (.A(G1757_490_gat), .B(G1794_460_gat), .Y(G2131_746_gat) );
AND2XL U_g698 (.A(G1764_488_gat), .B(G1794_460_gat), .Y(G2184_747_gat) );
AND2XL U_g699 (.A(G1771_485_gat), .B(G1794_460_gat), .Y(G2236_748_gat) );
AND2XL U_g700 (.A(G1495_672_gat), .B(G329_45_gat), .Y(G1503_749_gat) );
AND2XL U_g701 (.A(G1502_656_gat), .B(G326_44_gat), .Y(G1510_750_gat) );
AND2XL U_g702 (.A(G1478_671_gat), .B(G326_44_gat), .Y(G1486_751_gat) );
AND2XL U_g703 (.A(G1501_640_gat), .B(G322_43_gat), .Y(G1509_752_gat) );
AND2XL U_g704 (.A(G1485_655_gat), .B(G322_43_gat), .Y(G1493_753_gat) );
AND2XL U_g705 (.A(G1461_670_gat), .B(G322_43_gat), .Y(G1469_754_gat) );
AND2XL U_g706 (.A(G1500_720_gat), .B(G317_42_gat), .Y(G1508_755_gat) );
AND2XL U_g707 (.A(G1484_639_gat), .B(G317_42_gat), .Y(G1492_756_gat) );
AND2XL U_g708 (.A(G1468_654_gat), .B(G317_42_gat), .Y(G1476_757_gat) );
AND2XL U_g709 (.A(G1444_669_gat), .B(G317_42_gat), .Y(G1452_758_gat) );
AND2XL U_g710 (.A(G1499_704_gat), .B(G311_41_gat), .Y(G1507_759_gat) );
AND2XL U_g711 (.A(G1483_719_gat), .B(G311_41_gat), .Y(G1491_760_gat) );
AND2XL U_g712 (.A(G1467_638_gat), .B(G311_41_gat), .Y(G1475_761_gat) );
AND2XL U_g713 (.A(G1451_653_gat), .B(G311_41_gat), .Y(G1459_762_gat) );
AND2XL U_g714 (.A(G1427_668_gat), .B(G311_41_gat), .Y(G1435_763_gat) );
AND2XL U_g715 (.A(G1498_624_gat), .B(G303_40_gat), .Y(G1506_764_gat) );
AND2XL U_g716 (.A(G1482_703_gat), .B(G303_40_gat), .Y(G1490_765_gat) );
AND2XL U_g717 (.A(G1466_718_gat), .B(G303_40_gat), .Y(G1474_766_gat) );
AND2XL U_g718 (.A(G1450_637_gat), .B(G303_40_gat), .Y(G1458_767_gat) );
AND2XL U_g719 (.A(G1434_652_gat), .B(G303_40_gat), .Y(G1442_768_gat) );
AND2XL U_g720 (.A(G1410_667_gat), .B(G303_40_gat), .Y(G1418_769_gat) );
AND2XL U_g721 (.A(G1497_608_gat), .B(G294_39_gat), .Y(G1505_770_gat) );
AND2XL U_g722 (.A(G1481_623_gat), .B(G294_39_gat), .Y(G1489_771_gat) );
AND2XL U_g723 (.A(G1465_702_gat), .B(G294_39_gat), .Y(G1473_772_gat) );
AND2XL U_g724 (.A(G1449_717_gat), .B(G294_39_gat), .Y(G1457_773_gat) );
AND2XL U_g725 (.A(G1433_636_gat), .B(G294_39_gat), .Y(G1441_774_gat) );
AND2XL U_g726 (.A(G1417_651_gat), .B(G294_39_gat), .Y(G1425_775_gat) );
AND2XL U_g727 (.A(G1393_666_gat), .B(G294_39_gat), .Y(G1401_776_gat) );
AND2XL U_g728 (.A(G1496_688_gat), .B(G283_38_gat), .Y(G1504_777_gat) );
AND2XL U_g729 (.A(G1480_607_gat), .B(G283_38_gat), .Y(G1488_778_gat) );
AND2XL U_g730 (.A(G1464_622_gat), .B(G283_38_gat), .Y(G1472_779_gat) );
AND2XL U_g731 (.A(G1448_701_gat), .B(G283_38_gat), .Y(G1456_780_gat) );
AND2XL U_g732 (.A(G1432_716_gat), .B(G283_38_gat), .Y(G1440_781_gat) );
AND2XL U_g733 (.A(G1416_635_gat), .B(G283_38_gat), .Y(G1424_782_gat) );
AND2XL U_g734 (.A(G1400_650_gat), .B(G283_38_gat), .Y(G1408_783_gat) );
AND2XL U_g735 (.A(G1376_665_gat), .B(G283_38_gat), .Y(G1384_784_gat) );
AND3XL U_g736 (.A(G2236_748_ngat), .B(G2235_472_ngat), .C(G2234_480_ngat), .Y(G2237_785_gat) );
AND3XL U_g737 (.A(G2184_747_ngat), .B(G2183_473_ngat), .C(G2182_483_ngat), .Y(G2185_786_gat) );
AND3XL U_g738 (.A(G2131_746_ngat), .B(G2130_474_ngat), .C(G2129_484_ngat), .Y(G2132_787_gat) );
AND3XL U_g739 (.A(G2079_745_ngat), .B(G2078_475_ngat), .C(G2077_487_ngat), .Y(G2080_788_gat) );
AND3XL U_g740 (.A(G2024_744_ngat), .B(G2023_476_ngat), .C(G2022_489_ngat), .Y(G2025_789_gat) );
AND3XL U_g741 (.A(G1974_743_ngat), .B(G1973_477_ngat), .C(G1972_493_ngat), .Y(G1975_790_gat) );
AND3XL U_g742 (.A(G1923_742_ngat), .B(G1922_478_ngat), .C(G1921_495_ngat), .Y(G1924_791_gat) );
AND3XL U_g743 (.A(G1873_741_ngat), .B(G1872_479_ngat), .C(G1871_499_ngat), .Y(G1874_792_gat) );
AND2XL U_g744 (.A(G575_586_gat), .B(G574_585_gat), .Y(G576_793_gat) );
BUFX20 U_g745 (.A(G1029_588_gat), .Y(G360_794_gat) );
AND2XL U_g746 (.A(G2973_591_gat), .B(G2970_491_gat), .Y(G565_795_gat) );
AND2XL U_g747 (.A(G2981_592_gat), .B(G2978_492_gat), .Y(G569_796_gat) );
AND2XL U_g748 (.A(G2974_589_gat), .B(G2967_497_gat), .Y(G566_797_gat) );
AND2XL U_g749 (.A(G2982_590_gat), .B(G2975_498_gat), .Y(G570_798_gat) );
AND2XL U_g750 (.A(G1359_664_gat), .B(G159_21_gat), .Y(G1367_799_gat) );
AND2XL U_g751 (.A(G1349_647_gat), .B(G159_21_gat), .Y(G1357_800_gat) );
AND2XL U_g752 (.A(G1331_630_gat), .B(G159_21_gat), .Y(G1339_801_gat) );
AND2XL U_g753 (.A(G1313_709_gat), .B(G159_21_gat), .Y(G1321_802_gat) );
AND2XL U_g754 (.A(G1295_692_gat), .B(G159_21_gat), .Y(G1303_803_gat) );
AND2XL U_g755 (.A(G1277_611_gat), .B(G159_21_gat), .Y(G1285_804_gat) );
AND2XL U_g756 (.A(G1259_594_gat), .B(G159_21_gat), .Y(G1267_805_gat) );
AND2XL U_g757 (.A(G1241_673_gat), .B(G159_21_gat), .Y(G1249_806_gat) );
AND2XL U_g758 (.A(G1342_663_gat), .B(G150_20_gat), .Y(G1350_807_gat) );
AND2XL U_g759 (.A(G1332_646_gat), .B(G150_20_gat), .Y(G1340_808_gat) );
AND2XL U_g760 (.A(G1314_629_gat), .B(G150_20_gat), .Y(G1322_809_gat) );
AND2XL U_g761 (.A(G1296_708_gat), .B(G150_20_gat), .Y(G1304_810_gat) );
AND2XL U_g762 (.A(G1278_691_gat), .B(G150_20_gat), .Y(G1286_811_gat) );
AND2XL U_g763 (.A(G1260_610_gat), .B(G150_20_gat), .Y(G1268_812_gat) );
AND2XL U_g764 (.A(G1242_593_gat), .B(G150_20_gat), .Y(G1250_813_gat) );
AND2XL U_g765 (.A(G1325_662_gat), .B(G143_19_gat), .Y(G1333_814_gat) );
AND2XL U_g766 (.A(G1315_645_gat), .B(G143_19_gat), .Y(G1323_815_gat) );
AND2XL U_g767 (.A(G1297_628_gat), .B(G143_19_gat), .Y(G1305_816_gat) );
AND2XL U_g768 (.A(G1279_707_gat), .B(G143_19_gat), .Y(G1287_817_gat) );
AND2XL U_g769 (.A(G1261_690_gat), .B(G143_19_gat), .Y(G1269_818_gat) );
AND2XL U_g770 (.A(G1243_609_gat), .B(G143_19_gat), .Y(G1251_819_gat) );
AND2XL U_g771 (.A(G1308_661_gat), .B(G137_18_gat), .Y(G1316_820_gat) );
AND2XL U_g772 (.A(G1298_644_gat), .B(G137_18_gat), .Y(G1306_821_gat) );
AND2XL U_g773 (.A(G1280_627_gat), .B(G137_18_gat), .Y(G1288_822_gat) );
AND2XL U_g774 (.A(G1262_706_gat), .B(G137_18_gat), .Y(G1270_823_gat) );
AND2XL U_g775 (.A(G1244_689_gat), .B(G137_18_gat), .Y(G1252_824_gat) );
AND2XL U_g776 (.A(G1291_660_gat), .B(G132_17_gat), .Y(G1299_825_gat) );
AND2XL U_g777 (.A(G1281_643_gat), .B(G132_17_gat), .Y(G1289_826_gat) );
AND2XL U_g778 (.A(G1263_626_gat), .B(G132_17_gat), .Y(G1271_827_gat) );
AND2XL U_g779 (.A(G1245_705_gat), .B(G132_17_gat), .Y(G1253_828_gat) );
AND2XL U_g780 (.A(G1274_659_gat), .B(G128_16_gat), .Y(G1282_829_gat) );
AND2XL U_g781 (.A(G1264_642_gat), .B(G128_16_gat), .Y(G1272_830_gat) );
AND2XL U_g782 (.A(G1246_625_gat), .B(G128_16_gat), .Y(G1254_831_gat) );
AND2XL U_g783 (.A(G1257_658_gat), .B(G125_15_gat), .Y(G1265_832_gat) );
AND2XL U_g784 (.A(G1247_641_gat), .B(G125_15_gat), .Y(G1255_833_gat) );
AND2XL U_g785 (.A(G1240_657_gat), .B(G124_14_gat), .Y(G1248_834_gat) );
AND3XL U_g786 (.A(G2222_520_ngat), .B(G2219_380_ngat), .C(G2216_740_ngat), .Y(G2225_835_gat) );
AND3XL U_g787 (.A(G2222_520_ngat), .B(G2219_380_ngat), .C(G2216_740_ngat), .Y(G2229_836_gat) );
AND2XL U_g788 (.A(G3061_725_gat), .B(G3058_522_gat), .Y(G595_837_gat) );
AND2XL U_g789 (.A(G1383_649_gat), .B(G530_66_gat), .Y(G1391_838_gat) );
AND2XL U_g790 (.A(G1399_634_gat), .B(G530_66_gat), .Y(G1407_839_gat) );
AND2XL U_g791 (.A(G1415_715_gat), .B(G530_66_gat), .Y(G1423_840_gat) );
AND2XL U_g792 (.A(G1431_700_gat), .B(G530_66_gat), .Y(G1439_841_gat) );
AND2XL U_g793 (.A(G1447_621_gat), .B(G530_66_gat), .Y(G1455_842_gat) );
AND2XL U_g794 (.A(G1463_606_gat), .B(G530_66_gat), .Y(G1471_843_gat) );
AND2XL U_g795 (.A(G1479_687_gat), .B(G530_66_gat), .Y(G1487_844_gat) );
AND3XL U_g796 (.A(G2170_525_ngat), .B(G2167_384_ngat), .C(G2164_739_ngat), .Y(G2173_845_gat) );
AND3XL U_g797 (.A(G2170_525_ngat), .B(G2167_384_ngat), .C(G2164_739_ngat), .Y(G2177_846_gat) );
AND2XL U_g798 (.A(G1360_680_gat), .B(G517_70_gat), .Y(G1368_847_gat) );
AND2XL U_g799 (.A(G1382_633_gat), .B(G517_70_gat), .Y(G1390_848_gat) );
AND2XL U_g800 (.A(G1398_714_gat), .B(G517_70_gat), .Y(G1406_849_gat) );
AND2XL U_g801 (.A(G1414_699_gat), .B(G517_70_gat), .Y(G1422_850_gat) );
AND2XL U_g802 (.A(G1430_620_gat), .B(G517_70_gat), .Y(G1438_851_gat) );
AND2XL U_g803 (.A(G1446_605_gat), .B(G517_70_gat), .Y(G1454_852_gat) );
AND2XL U_g804 (.A(G1462_686_gat), .B(G517_70_gat), .Y(G1470_853_gat) );
AND2XL U_g805 (.A(G3062_721_gat), .B(G3055_532_gat), .Y(G596_854_gat) );
AND2XL U_g806 (.A(G1343_679_gat), .B(G504_76_gat), .Y(G1351_855_gat) );
AND2XL U_g807 (.A(G1361_600_gat), .B(G504_76_gat), .Y(G1369_856_gat) );
AND2XL U_g808 (.A(G1381_713_gat), .B(G504_76_gat), .Y(G1389_857_gat) );
AND2XL U_g809 (.A(G1397_698_gat), .B(G504_76_gat), .Y(G1405_858_gat) );
AND2XL U_g810 (.A(G1413_619_gat), .B(G504_76_gat), .Y(G1421_859_gat) );
AND2XL U_g811 (.A(G1429_604_gat), .B(G504_76_gat), .Y(G1437_860_gat) );
AND2XL U_g812 (.A(G1445_685_gat), .B(G504_76_gat), .Y(G1453_861_gat) );
AND3XL U_g813 (.A(G2065_534_ngat), .B(G2062_395_ngat), .C(G2059_738_ngat), .Y(G2068_862_gat) );
AND3XL U_g814 (.A(G2065_534_ngat), .B(G2062_395_ngat), .C(G2059_738_ngat), .Y(G2072_863_gat) );
AND2XL U_g815 (.A(G1326_678_gat), .B(G492_80_gat), .Y(G1334_864_gat) );
AND2XL U_g816 (.A(G1344_599_gat), .B(G492_80_gat), .Y(G1352_865_gat) );
AND2XL U_g817 (.A(G1362_616_gat), .B(G492_80_gat), .Y(G1370_866_gat) );
AND2XL U_g818 (.A(G1380_697_gat), .B(G492_80_gat), .Y(G1388_867_gat) );
AND2XL U_g819 (.A(G1396_618_gat), .B(G492_80_gat), .Y(G1404_868_gat) );
AND2XL U_g820 (.A(G1412_603_gat), .B(G492_80_gat), .Y(G1420_869_gat) );
AND2XL U_g821 (.A(G1428_684_gat), .B(G492_80_gat), .Y(G1436_870_gat) );
AND3XL U_g822 (.A(G2010_537_ngat), .B(G2007_401_ngat), .C(G2004_737_ngat), .Y(G2013_871_gat) );
AND3XL U_g823 (.A(G2010_537_ngat), .B(G2007_401_ngat), .C(G2004_737_ngat), .Y(G2017_872_gat) );
AND2XL U_g824 (.A(G1309_677_gat), .B(G483_81_gat), .Y(G1317_873_gat) );
AND2XL U_g825 (.A(G1327_598_gat), .B(G483_81_gat), .Y(G1335_874_gat) );
AND2XL U_g826 (.A(G1345_615_gat), .B(G483_81_gat), .Y(G1353_875_gat) );
AND2XL U_g827 (.A(G1363_696_gat), .B(G483_81_gat), .Y(G1371_876_gat) );
AND2XL U_g828 (.A(G1379_617_gat), .B(G483_81_gat), .Y(G1387_877_gat) );
AND2XL U_g829 (.A(G1395_602_gat), .B(G483_81_gat), .Y(G1403_878_gat) );
AND2XL U_g830 (.A(G1411_683_gat), .B(G483_81_gat), .Y(G1419_879_gat) );
AND2XL U_g831 (.A(G3053_731_gat), .B(G3050_539_gat), .Y(G589_880_gat) );
AND3XL U_g832 (.A(G1960_540_ngat), .B(G1957_407_ngat), .C(G1954_736_ngat), .Y(G1963_881_gat) );
AND3XL U_g833 (.A(G1960_540_ngat), .B(G1957_407_ngat), .C(G1954_736_ngat), .Y(G1967_882_gat) );
AND2XL U_g834 (.A(G1292_676_gat), .B(G467_87_gat), .Y(G1300_883_gat) );
AND2XL U_g835 (.A(G1310_597_gat), .B(G467_87_gat), .Y(G1318_884_gat) );
AND2XL U_g836 (.A(G1328_614_gat), .B(G467_87_gat), .Y(G1336_885_gat) );
AND2XL U_g837 (.A(G1346_695_gat), .B(G467_87_gat), .Y(G1354_886_gat) );
AND2XL U_g838 (.A(G1364_712_gat), .B(G467_87_gat), .Y(G1372_887_gat) );
AND2XL U_g839 (.A(G1378_601_gat), .B(G467_87_gat), .Y(G1386_888_gat) );
AND2XL U_g840 (.A(G1394_682_gat), .B(G467_87_gat), .Y(G1402_889_gat) );
AND2XL U_g841 (.A(G644_269_ngat), .B(G641_728_ngat), .Y(G645_890_gat) );
AND2XL U_g842 (.A(G3054_726_gat), .B(G3047_546_gat), .Y(G590_891_gat) );
AND2XL U_g843 (.A(G1275_675_gat), .B(G447_95_gat), .Y(G1283_892_gat) );
AND2XL U_g844 (.A(G1293_596_gat), .B(G447_95_gat), .Y(G1301_893_gat) );
AND2XL U_g845 (.A(G1311_613_gat), .B(G447_95_gat), .Y(G1319_894_gat) );
AND2XL U_g846 (.A(G1329_694_gat), .B(G447_95_gat), .Y(G1337_895_gat) );
AND2XL U_g847 (.A(G1347_711_gat), .B(G447_95_gat), .Y(G1355_896_gat) );
AND2XL U_g848 (.A(G1365_632_gat), .B(G447_95_gat), .Y(G1373_897_gat) );
AND2XL U_g849 (.A(G1377_681_gat), .B(G447_95_gat), .Y(G1385_898_gat) );
AND3XL U_g850 (.A(G1859_547_ngat), .B(G1856_417_ngat), .C(G1853_735_ngat), .Y(G1862_899_gat) );
AND3XL U_g851 (.A(G1859_547_ngat), .B(G1856_417_ngat), .C(G1853_735_ngat), .Y(G1866_900_gat) );
AND2XL U_g852 (.A(G1258_674_gat), .B(G432_99_gat), .Y(G1266_901_gat) );
AND2XL U_g853 (.A(G1276_595_gat), .B(G432_99_gat), .Y(G1284_902_gat) );
AND2XL U_g854 (.A(G1294_612_gat), .B(G432_99_gat), .Y(G1302_903_gat) );
AND2XL U_g855 (.A(G1312_693_gat), .B(G432_99_gat), .Y(G1320_904_gat) );
AND2XL U_g856 (.A(G1330_710_gat), .B(G432_99_gat), .Y(G1338_905_gat) );
AND2XL U_g857 (.A(G1348_631_gat), .B(G432_99_gat), .Y(G1356_906_gat) );
AND2XL U_g858 (.A(G1366_648_gat), .B(G432_99_gat), .Y(G1374_907_gat) );
AND2XL U_g859 (.A(G980_200_gat), .B(G902_729_gat), .Y(G983_908_gat) );
AND2XL U_g860 (.A(G1008_204_gat), .B(G911_724_gat), .Y(G1011_909_gat) );
AND2XL U_g861 (.A(G942_441_gat), .B(G649_723_gat), .Y(G947_910_gat) );
AND8XL U_g862 (.A(G1510_750_ngat), .B(G1509_752_ngat), .C(G1508_755_ngat), .D(G1507_759_ngat), .E(G1506_764_ngat), .F(G1505_770_ngat), .G(G1504_777_ngat), .H(G1503_749_ngat), .Y(G1511_911_gat) );
AND8XL U_g863 (.A(G1493_753_ngat), .B(G1492_756_ngat), .C(G1491_760_ngat), .D(G1490_765_ngat), .E(G1489_771_ngat), .F(G1488_778_ngat), .G(G1487_844_ngat), .H(G1486_751_ngat), .Y(G1494_912_gat) );
AND8XL U_g864 (.A(G1476_757_ngat), .B(G1475_761_ngat), .C(G1474_766_ngat), .D(G1473_772_ngat), .E(G1472_779_ngat), .F(G1471_843_ngat), .G(G1470_853_ngat), .H(G1469_754_ngat), .Y(G1477_913_gat) );
AND8XL U_g865 (.A(G1459_762_ngat), .B(G1458_767_ngat), .C(G1457_773_ngat), .D(G1456_780_ngat), .E(G1455_842_ngat), .F(G1454_852_ngat), .G(G1453_861_ngat), .H(G1452_758_ngat), .Y(G1460_914_gat) );
AND8XL U_g866 (.A(G1442_768_ngat), .B(G1441_774_ngat), .C(G1440_781_ngat), .D(G1439_841_ngat), .E(G1438_851_ngat), .F(G1437_860_ngat), .G(G1436_870_ngat), .H(G1435_763_ngat), .Y(G1443_915_gat) );
AND8XL U_g867 (.A(G1425_775_ngat), .B(G1424_782_ngat), .C(G1423_840_ngat), .D(G1422_850_ngat), .E(G1421_859_ngat), .F(G1420_869_ngat), .G(G1419_879_ngat), .H(G1418_769_ngat), .Y(G1426_916_gat) );
AND8XL U_g868 (.A(G1408_783_ngat), .B(G1407_839_ngat), .C(G1406_849_ngat), .D(G1405_858_ngat), .E(G1404_868_ngat), .F(G1403_878_ngat), .G(G1402_889_ngat), .H(G1401_776_ngat), .Y(G1409_917_gat) );
AND8XL U_g869 (.A(G1391_838_ngat), .B(G1390_848_ngat), .C(G1389_857_ngat), .D(G1388_867_ngat), .E(G1387_877_ngat), .F(G1386_888_ngat), .G(G1385_898_ngat), .H(G1384_784_ngat), .Y(G1392_918_gat) );
BUFX20 U_g870 (.A(G2237_785_gat), .Y(G2242_919_gat) );
BUFX20 U_g871 (.A(G2237_785_gat), .Y(G2245_920_gat) );
BUFX20 U_g872 (.A(G2237_785_gat), .Y(G2477_921_gat) );
BUFX20 U_g873 (.A(G2185_786_gat), .Y(G2190_922_gat) );
BUFX20 U_g874 (.A(G2185_786_gat), .Y(G2193_923_gat) );
BUFX20 U_g875 (.A(G2185_786_gat), .Y(G2476_924_gat) );
BUFX20 U_g876 (.A(G2132_787_gat), .Y(G2137_925_gat) );
BUFX20 U_g877 (.A(G2132_787_gat), .Y(G2140_926_gat) );
BUFX20 U_g878 (.A(G2132_787_gat), .Y(G2475_927_gat) );
BUFX20 U_g879 (.A(G2080_788_gat), .Y(G2085_928_gat) );
BUFX20 U_g880 (.A(G2080_788_gat), .Y(G2088_929_gat) );
BUFX20 U_g881 (.A(G2080_788_gat), .Y(G2474_930_gat) );
BUFX20 U_g882 (.A(G2025_789_gat), .Y(G2028_931_gat) );
BUFX20 U_g883 (.A(G2025_789_gat), .Y(G2031_932_gat) );
BUFX20 U_g884 (.A(G1975_790_gat), .Y(G1978_933_gat) );
BUFX20 U_g885 (.A(G1975_790_gat), .Y(G1981_934_gat) );
BUFX20 U_g886 (.A(G1924_791_gat), .Y(G1927_935_gat) );
BUFX20 U_g887 (.A(G1924_791_gat), .Y(G1930_936_gat) );
BUFX20 U_g888 (.A(G1874_792_gat), .Y(G1877_937_gat) );
BUFX20 U_g889 (.A(G1874_792_gat), .Y(G1880_938_gat) );
BUFX20 U_g890 (.A(G576_793_gat), .Y(G579_939_gat) );
AND2XL U_g891 (.A(G360_794_gat), .B(G359_587_gat), .Y(G361_940_gat) );
AND2XL U_g892 (.A(G566_797_gat), .B(G565_795_gat), .Y(G567_941_gat) );
AND2XL U_g893 (.A(G570_798_gat), .B(G569_796_gat), .Y(G571_942_gat) );
AND2XL U_g894 (.A(G2173_845_gat), .B(G2298_237_gat), .Y(G2383_943_gat) );
AND2XL U_g895 (.A(G2225_835_gat), .B(G2298_237_gat), .Y(G2391_944_gat) );
AND2XL U_g896 (.A(G1963_881_gat), .B(G2289_239_gat), .Y(G2341_945_gat) );
AND2XL U_g897 (.A(G2013_871_gat), .B(G2289_239_gat), .Y(G2354_946_gat) );
AND2XL U_g898 (.A(G2068_862_gat), .B(G2289_239_gat), .Y(G2367_947_gat) );
AND2XL U_g899 (.A(G1862_899_gat), .B(G2285_241_gat), .Y(G2320_948_gat) );
AND5XL U_g900 (.A(G2481_150_gat), .B(G2237_785_gat), .C(G2185_786_gat), .D(G2132_787_gat), .E(G2080_788_gat), .Y(G2482_949_gat) );
AND8XL U_g901 (.A(G1374_907_ngat), .B(G1373_897_ngat), .C(G1372_887_ngat), .D(G1371_876_ngat), .E(G1370_866_ngat), .F(G1369_856_ngat), .G(G1368_847_ngat), .H(G1367_799_ngat), .Y(G1375_950_gat) );
AND8XL U_g902 (.A(G1357_800_ngat), .B(G1356_906_ngat), .C(G1355_896_ngat), .D(G1354_886_ngat), .E(G1353_875_ngat), .F(G1352_865_ngat), .G(G1351_855_ngat), .H(G1350_807_ngat), .Y(G1358_951_gat) );
AND8XL U_g903 (.A(G1340_808_ngat), .B(G1339_801_ngat), .C(G1338_905_ngat), .D(G1337_895_ngat), .E(G1336_885_ngat), .F(G1335_874_ngat), .G(G1334_864_ngat), .H(G1333_814_ngat), .Y(G1341_952_gat) );
AND8XL U_g904 (.A(G1323_815_ngat), .B(G1322_809_ngat), .C(G1321_802_ngat), .D(G1320_904_ngat), .E(G1319_894_ngat), .F(G1318_884_ngat), .G(G1317_873_ngat), .H(G1316_820_ngat), .Y(G1324_953_gat) );
AND8XL U_g905 (.A(G1306_821_ngat), .B(G1305_816_ngat), .C(G1304_810_ngat), .D(G1303_803_ngat), .E(G1302_903_ngat), .F(G1301_893_ngat), .G(G1300_883_ngat), .H(G1299_825_ngat), .Y(G1307_954_gat) );
AND8XL U_g906 (.A(G1289_826_ngat), .B(G1288_822_ngat), .C(G1287_817_ngat), .D(G1286_811_ngat), .E(G1285_804_ngat), .F(G1284_902_ngat), .G(G1283_892_ngat), .H(G1282_829_ngat), .Y(G1290_955_gat) );
AND8XL U_g907 (.A(G1272_830_ngat), .B(G1271_827_ngat), .C(G1270_823_ngat), .D(G1269_818_ngat), .E(G1268_812_ngat), .F(G1267_805_ngat), .G(G1266_901_ngat), .H(G1265_832_ngat), .Y(G1273_956_gat) );
AND8XL U_g908 (.A(G1255_833_ngat), .B(G1254_831_ngat), .C(G1253_828_ngat), .D(G1252_824_ngat), .E(G1251_819_ngat), .F(G1250_813_ngat), .G(G1249_806_ngat), .H(G1248_834_ngat), .Y(G1256_957_gat) );
AND3XL U_g909 (.A(G985_378_ngat), .B(G984_408_ngat), .C(G983_908_ngat), .Y(G986_958_gat) );
BUFX20 U_g910 (.A(G2229_836_gat), .Y(G2256_959_gat) );
AND2XL U_g911 (.A(G596_854_gat), .B(G595_837_gat), .Y(G597_960_gat) );
BUFX20 U_g912 (.A(G2177_846_gat), .Y(G2204_961_gat) );
AND3XL U_g913 (.A(G1013_403_ngat), .B(G1012_386_ngat), .C(G1011_909_ngat), .Y(G1014_962_gat) );
BUFX20 U_g914 (.A(G2072_863_gat), .Y(G2099_963_gat) );
BUFX20 U_g915 (.A(G2017_872_gat), .Y(G2042_964_gat) );
AND2XL U_g916 (.A(G590_891_gat), .B(G589_880_gat), .Y(G591_965_gat) );
BUFX20 U_g917 (.A(G1967_882_gat), .Y(G1992_966_gat) );
BUFX20 U_g918 (.A(G1866_900_gat), .Y(G1891_967_gat) );
AND2XL U_g919 (.A(G610_432_gat), .B(G576_793_gat), .Y(G614_968_gat) );
AND2XL U_g920 (.A(G941_333_gat), .B(G645_890_gat), .Y(G944_969_gat) );
BUFX20 U_g921 (.A(G579_939_gat), .Y(G2994_970_gat) );
BUFX20 U_g922 (.A(G579_939_gat), .Y(G3002_971_gat) );
BUFX20 U_g923 (.A(G567_941_gat), .Y(G568_972_gat) );
BUFX20 U_g924 (.A(G571_942_gat), .Y(G2991_973_gat) );
BUFX20 U_g925 (.A(G571_942_gat), .Y(G2999_974_gat) );
BUFX20 U_g926 (.A(G2383_943_gat), .Y(G3224_975_gat) );
BUFX20 U_g927 (.A(G2383_943_gat), .Y(G3232_976_gat) );
BUFX20 U_g928 (.A(G2391_944_gat), .Y(G3240_977_gat) );
BUFX20 U_g929 (.A(G2391_944_gat), .Y(G3248_978_gat) );
BUFX20 U_g930 (.A(G2341_945_gat), .Y(G3158_979_gat) );
BUFX20 U_g931 (.A(G2341_945_gat), .Y(G3166_980_gat) );
BUFX20 U_g932 (.A(G2354_946_gat), .Y(G3174_981_gat) );
BUFX20 U_g933 (.A(G2354_946_gat), .Y(G3182_982_gat) );
BUFX20 U_g934 (.A(G2367_947_gat), .Y(G3190_983_gat) );
BUFX20 U_g935 (.A(G2367_947_gat), .Y(G3200_984_gat) );
BUFX20 U_g936 (.A(G2320_948_gat), .Y(G3124_985_gat) );
BUFX20 U_g937 (.A(G2320_948_gat), .Y(G3134_986_gat) );
AND3XL U_g938 (.A(G2242_919_gat), .B(G2229_836_gat), .C(G200_25_gat), .Y(G2255_987_gat) );
AND3XL U_g939 (.A(G2190_922_gat), .B(G2177_846_gat), .C(G200_25_gat), .Y(G2203_988_gat) );
AND3XL U_g940 (.A(G2085_928_gat), .B(G2072_863_gat), .C(G200_25_gat), .Y(G2098_989_gat) );
AND3XL U_g941 (.A(G2028_931_gat), .B(G2017_872_gat), .C(G200_25_gat), .Y(G2041_990_gat) );
AND3XL U_g942 (.A(G1978_933_gat), .B(G1967_882_gat), .C(G200_25_gat), .Y(G1991_991_gat) );
AND3XL U_g943 (.A(G1877_937_gat), .B(G1866_900_gat), .C(G200_25_gat), .Y(G1890_992_gat) );
AND3XL U_g944 (.A(G2245_920_gat), .B(G2229_836_gat), .C(G190_24_gat), .Y(G2254_993_gat) );
AND3XL U_g945 (.A(G2193_923_gat), .B(G2177_846_gat), .C(G190_24_gat), .Y(G2202_994_gat) );
AND3XL U_g946 (.A(G2088_929_gat), .B(G2072_863_gat), .C(G190_24_gat), .Y(G2097_995_gat) );
AND3XL U_g947 (.A(G2031_932_gat), .B(G2017_872_gat), .C(G190_24_gat), .Y(G2040_996_gat) );
AND3XL U_g948 (.A(G1981_934_gat), .B(G1967_882_gat), .C(G190_24_gat), .Y(G1990_997_gat) );
AND3XL U_g949 (.A(G1880_938_gat), .B(G1866_900_gat), .C(G190_24_gat), .Y(G1889_998_gat) );
AND5XL U_g950 (.A(G2478_64_gat), .B(G2477_921_gat), .C(G2476_924_gat), .D(G2475_927_gat), .E(G2474_930_gat), .Y(G2483_999_gat) );
AND3XL U_g951 (.A(G2245_920_gat), .B(G2225_835_gat), .C(G179_23_gat), .Y(G2251_1000_gat) );
AND3XL U_g952 (.A(G2193_923_gat), .B(G2173_845_gat), .C(G179_23_gat), .Y(G2199_1001_gat) );
AND3XL U_g953 (.A(G2088_929_gat), .B(G2068_862_gat), .C(G179_23_gat), .Y(G2094_1002_gat) );
AND3XL U_g954 (.A(G2031_932_gat), .B(G2013_871_gat), .C(G179_23_gat), .Y(G2037_1003_gat) );
AND3XL U_g955 (.A(G1981_934_gat), .B(G1963_881_gat), .C(G179_23_gat), .Y(G1987_1004_gat) );
AND3XL U_g956 (.A(G1880_938_gat), .B(G1862_899_gat), .C(G179_23_gat), .Y(G1886_1005_gat) );
AND3XL U_g957 (.A(G2242_919_gat), .B(G2225_835_gat), .C(G169_22_gat), .Y(G2248_1006_gat) );
AND3XL U_g958 (.A(G2190_922_gat), .B(G2173_845_gat), .C(G169_22_gat), .Y(G2196_1007_gat) );
AND3XL U_g959 (.A(G2085_928_gat), .B(G2068_862_gat), .C(G169_22_gat), .Y(G2091_1008_gat) );
AND3XL U_g960 (.A(G2028_931_gat), .B(G2013_871_gat), .C(G169_22_gat), .Y(G2034_1009_gat) );
AND3XL U_g961 (.A(G1978_933_gat), .B(G1963_881_gat), .C(G169_22_gat), .Y(G1984_1010_gat) );
AND3XL U_g962 (.A(G1877_937_gat), .B(G1862_899_gat), .C(G169_22_gat), .Y(G1883_1011_gat) );
BUFX20 U_g963 (.A(G597_960_gat), .Y(G600_1012_gat) );
BUFX20 U_g964 (.A(G591_965_gat), .Y(G3063_1013_gat) );
BUFX20 U_g965 (.A(G591_965_gat), .Y(G3071_1014_gat) );
AND2XL U_g966 (.A(G678_275_gat), .B(G591_965_gat), .Y(G679_1015_gat) );
AND2XL U_g967 (.A(G1533_421_gat), .B(G1256_957_gat), .Y(G1536_1016_gat) );
AND3XL U_g968 (.A(G617_536_ngat), .B(G616_424_ngat), .C(G614_968_ngat), .Y(G618_1017_gat) );
AND2XL U_g969 (.A(G1534_431_gat), .B(G1392_918_gat), .Y(G1537_1018_gat) );
AND2XL U_g970 (.A(G665_433_gat), .B(G597_960_gat), .Y(G669_1019_gat) );
AND2XL U_g971 (.A(G1581_304_gat), .B(G1273_956_gat), .Y(G1582_1020_gat) );
AND2XL U_g972 (.A(G1512_193_gat), .B(G1409_917_gat), .Y(G1583_1021_gat) );
AND2XL U_g973 (.A(G1585_305_gat), .B(G1290_955_gat), .Y(G1586_1022_gat) );
AND2XL U_g974 (.A(G1512_193_gat), .B(G1426_916_gat), .Y(G1587_1023_gat) );
AND2XL U_g975 (.A(G1589_306_gat), .B(G1307_954_gat), .Y(G1590_1024_gat) );
AND2XL U_g976 (.A(G1512_193_gat), .B(G1443_915_gat), .Y(G1591_1025_gat) );
AND2XL U_g977 (.A(G1593_307_gat), .B(G1324_953_gat), .Y(G1594_1026_gat) );
AND2XL U_g978 (.A(G1512_193_gat), .B(G1460_914_gat), .Y(G1595_1027_gat) );
AND2XL U_g979 (.A(G1597_308_gat), .B(G1341_952_gat), .Y(G1598_1028_gat) );
AND2XL U_g980 (.A(G1512_193_gat), .B(G1477_913_gat), .Y(G1599_1029_gat) );
AND2XL U_g981 (.A(G1601_309_gat), .B(G1358_951_gat), .Y(G1602_1030_gat) );
AND2XL U_g982 (.A(G1512_193_gat), .B(G1494_912_gat), .Y(G1603_1031_gat) );
AND2XL U_g983 (.A(G1605_310_gat), .B(G1375_950_gat), .Y(G1606_1032_gat) );
AND2XL U_g984 (.A(G1512_193_gat), .B(G1511_911_gat), .Y(G1607_1033_gat) );
AND2XL U_g985 (.A(G1901_336_gat), .B(G986_958_gat), .Y(G1903_1034_gat) );
AND2XL U_g986 (.A(G2109_340_gat), .B(G1014_962_gat), .Y(G2111_1035_gat) );
BUFX20 U_g987 (.A(G2994_970_gat), .Y(G2998_1036_gat) );
BUFX20 U_g988 (.A(G3002_971_gat), .Y(G3006_1037_gat) );
BUFX20 U_g989 (.A(G2991_973_gat), .Y(G2997_1038_gat) );
BUFX20 U_g990 (.A(G2999_974_gat), .Y(G3005_1039_gat) );
BUFX20 U_g991 (.A(G3224_975_gat), .Y(G3228_1040_gat) );
BUFX20 U_g992 (.A(G3232_976_gat), .Y(G3236_1041_gat) );
BUFX20 U_g993 (.A(G3240_977_gat), .Y(G3244_1042_gat) );
BUFX20 U_g994 (.A(G3248_978_gat), .Y(G3252_1043_gat) );
BUFX20 U_g995 (.A(G3158_979_gat), .Y(G3162_1044_gat) );
BUFX20 U_g996 (.A(G3166_980_gat), .Y(G3170_1045_gat) );
BUFX20 U_g997 (.A(G3174_981_gat), .Y(G3178_1046_gat) );
BUFX20 U_g998 (.A(G3182_982_gat), .Y(G3186_1047_gat) );
BUFX20 U_g999 (.A(G3190_983_gat), .Y(G3194_1048_gat) );
BUFX20 U_g1000 (.A(G3200_984_gat), .Y(G3204_1049_gat) );
BUFX20 U_g1001 (.A(G3124_985_gat), .Y(G3128_1050_gat) );
BUFX20 U_g1002 (.A(G3134_986_gat), .Y(G3138_1051_gat) );
AND2XL U_g1003 (.A(G2483_999_ngat), .B(G2482_949_ngat), .Y(G2484_1052_gat) );
AND2XL U_g1004 (.A(G2251_1000_ngat), .B(G2248_1006_ngat), .Y(G2257_1053_gat) );
AND2XL U_g1005 (.A(G2251_1000_ngat), .B(G2248_1006_ngat), .Y(G2260_1054_gat) );
AND2XL U_g1006 (.A(G2199_1001_ngat), .B(G2196_1007_ngat), .Y(G2205_1055_gat) );
AND2XL U_g1007 (.A(G2199_1001_ngat), .B(G2196_1007_ngat), .Y(G2208_1056_gat) );
AND2XL U_g1008 (.A(G2094_1002_ngat), .B(G2091_1008_ngat), .Y(G2100_1057_gat) );
AND2XL U_g1009 (.A(G2094_1002_ngat), .B(G2091_1008_ngat), .Y(G2101_1058_gat) );
AND2XL U_g1010 (.A(G2037_1003_ngat), .B(G2034_1009_ngat), .Y(G2043_1059_gat) );
AND2XL U_g1011 (.A(G2037_1003_ngat), .B(G2034_1009_ngat), .Y(G2046_1060_gat) );
AND2XL U_g1012 (.A(G1987_1004_ngat), .B(G1984_1010_ngat), .Y(G1993_1061_gat) );
AND2XL U_g1013 (.A(G1987_1004_ngat), .B(G1984_1010_ngat), .Y(G1996_1062_gat) );
AND2XL U_g1014 (.A(G1886_1005_ngat), .B(G1883_1011_ngat), .Y(G1892_1063_gat) );
AND2XL U_g1015 (.A(G1886_1005_ngat), .B(G1883_1011_ngat), .Y(G1893_1064_gat) );
AND3XL U_g1016 (.A(G2256_959_ngat), .B(G2255_987_ngat), .C(G2254_993_ngat), .Y(G2261_1065_gat) );
BUFX20 U_g1017 (.A(G600_1012_gat), .Y(G3066_1066_gat) );
BUFX20 U_g1018 (.A(G600_1012_gat), .Y(G3074_1067_gat) );
AND3XL U_g1019 (.A(G2204_961_ngat), .B(G2203_988_ngat), .C(G2202_994_ngat), .Y(G2209_1068_gat) );
AND3XL U_g1020 (.A(G2117_531_ngat), .B(G2114_388_ngat), .C(G2111_1035_ngat), .Y(G2120_1069_gat) );
AND3XL U_g1021 (.A(G2117_531_ngat), .B(G2114_388_ngat), .C(G2111_1035_ngat), .Y(G2124_1070_gat) );
AND3XL U_g1022 (.A(G2099_963_ngat), .B(G2098_989_ngat), .C(G2097_995_ngat), .Y(G2102_1071_gat) );
AND3XL U_g1023 (.A(G2042_964_ngat), .B(G2041_990_ngat), .C(G2040_996_ngat), .Y(G2047_1072_gat) );
BUFX20 U_g1024 (.A(G3063_1013_gat), .Y(G3069_1073_gat) );
BUFX20 U_g1025 (.A(G3071_1014_gat), .Y(G3077_1074_gat) );
AND3XL U_g1026 (.A(G1992_966_ngat), .B(G1991_991_ngat), .C(G1990_997_ngat), .Y(G1997_1075_gat) );
AND3XL U_g1027 (.A(G1909_545_ngat), .B(G1906_411_ngat), .C(G1903_1034_ngat), .Y(G1912_1076_gat) );
AND3XL U_g1028 (.A(G1909_545_ngat), .B(G1906_411_ngat), .C(G1903_1034_ngat), .Y(G1916_1077_gat) );
AND3XL U_g1029 (.A(G1891_967_ngat), .B(G1890_992_ngat), .C(G1889_998_ngat), .Y(G1894_1078_gat) );
AND3XL U_g1030 (.A(G1538_548_ngat), .B(G1537_1018_ngat), .C(G1536_1016_ngat), .Y(G1539_1079_gat) );
AND2XL U_g1031 (.A(G660_274_gat), .B(G568_972_gat), .Y(G661_1080_gat) );
AND2XL U_g1032 (.A(G680_420_ngat), .B(G679_1015_ngat), .Y(G681_1081_gat) );
AND3XL U_g1033 (.A(G672_533_ngat), .B(G671_426_ngat), .C(G669_1019_ngat), .Y(G673_1082_gat) );
AND2XL U_g1034 (.A(G1583_1021_ngat), .B(G1582_1020_ngat), .Y(G1584_1083_gat) );
AND2XL U_g1035 (.A(G1587_1023_ngat), .B(G1586_1022_ngat), .Y(G1588_1084_gat) );
AND2XL U_g1036 (.A(G1591_1025_ngat), .B(G1590_1024_ngat), .Y(G1592_1085_gat) );
AND2XL U_g1037 (.A(G1595_1027_ngat), .B(G1594_1026_ngat), .Y(G1596_1086_gat) );
AND2XL U_g1038 (.A(G1599_1029_ngat), .B(G1598_1028_ngat), .Y(G1600_1087_gat) );
AND2XL U_g1039 (.A(G1603_1031_ngat), .B(G1602_1030_ngat), .Y(G1604_1088_gat) );
AND2XL U_g1040 (.A(G1607_1033_ngat), .B(G1606_1032_ngat), .Y(G1608_1089_gat) );
AND2XL U_g1041 (.A(G1647_551_gat), .B(G618_1017_gat), .Y(G1652_1090_gat) );
AND2XL U_g1042 (.A(G2997_1038_gat), .B(G2994_970_gat), .Y(G619_1091_gat) );
AND2XL U_g1043 (.A(G3005_1039_gat), .B(G3002_971_gat), .Y(G582_1092_gat) );
AND2XL U_g1044 (.A(G2998_1036_gat), .B(G2991_973_gat), .Y(G620_1093_gat) );
AND2XL U_g1045 (.A(G3006_1037_gat), .B(G2999_974_gat), .Y(G583_1094_gat) );
AND2XL U_g1046 (.A(G2302_236_gat), .B(G2205_1055_gat), .Y(G2455_1095_gat) );
AND2XL U_g1047 (.A(G2302_236_gat), .B(G2257_1053_gat), .Y(G2458_1096_gat) );
AND2XL U_g1048 (.A(G2120_1069_gat), .B(G2298_237_gat), .Y(G2375_1097_gat) );
AND2XL U_g1049 (.A(G2293_238_gat), .B(G1993_1061_gat), .Y(G2445_1098_gat) );
AND2XL U_g1050 (.A(G2293_238_gat), .B(G2043_1059_gat), .Y(G2448_1099_gat) );
AND2XL U_g1051 (.A(G2488_503_gat), .B(G2484_1052_gat), .Y(G2489_1100_gat) );
AND2XL U_g1052 (.A(G1912_1076_gat), .B(G2285_241_gat), .Y(G2328_1101_gat) );
AND3XL U_g1053 (.A(G2137_925_gat), .B(G2124_1070_gat), .C(G200_25_gat), .Y(G2150_1102_gat) );
AND3XL U_g1054 (.A(G1927_935_gat), .B(G1916_1077_gat), .C(G200_25_gat), .Y(G1940_1103_gat) );
AND3XL U_g1055 (.A(G2140_926_gat), .B(G2124_1070_gat), .C(G190_24_gat), .Y(G2149_1104_gat) );
AND3XL U_g1056 (.A(G1930_936_gat), .B(G1916_1077_gat), .C(G190_24_gat), .Y(G1939_1105_gat) );
AND2XL U_g1057 (.A(G2261_1065_gat), .B(G2260_1054_gat), .Y(G2262_1106_gat) );
AND2XL U_g1058 (.A(G2209_1068_gat), .B(G2208_1056_gat), .Y(G2210_1107_gat) );
AND3XL U_g1059 (.A(G2140_926_gat), .B(G2120_1069_gat), .C(G179_23_gat), .Y(G2146_1108_gat) );
BUFX20 U_g1060 (.A(G2100_1057_gat), .Y(G2311_1109_gat) );
AND2XL U_g1061 (.A(G2102_1071_gat), .B(G2101_1058_gat), .Y(G2103_1110_gat) );
AND2XL U_g1062 (.A(G2047_1072_gat), .B(G2046_1060_gat), .Y(G2048_1111_gat) );
AND2XL U_g1063 (.A(G1997_1075_gat), .B(G1996_1062_gat), .Y(G1998_1112_gat) );
AND3XL U_g1064 (.A(G1930_936_gat), .B(G1912_1076_gat), .C(G179_23_gat), .Y(G1936_1113_gat) );
BUFX20 U_g1065 (.A(G1892_1063_gat), .Y(G2271_1114_gat) );
AND2XL U_g1066 (.A(G1894_1078_gat), .B(G1893_1064_gat), .Y(G1895_1115_gat) );
AND3XL U_g1067 (.A(G2137_925_gat), .B(G2120_1069_gat), .C(G169_22_gat), .Y(G2143_1116_gat) );
AND3XL U_g1068 (.A(G1927_935_gat), .B(G1912_1076_gat), .C(G169_22_gat), .Y(G1933_1117_gat) );
AND2XL U_g1069 (.A(G3069_1073_gat), .B(G3066_1066_gat), .Y(G606_1118_gat) );
BUFX20 U_g1070 (.A(G3066_1066_gat), .Y(G3070_1119_gat) );
AND2XL U_g1071 (.A(G3077_1074_gat), .B(G3074_1067_gat), .Y(G603_1120_gat) );
BUFX20 U_g1072 (.A(G3074_1067_gat), .Y(G3078_1121_gat) );
BUFX20 U_g1073 (.A(G2124_1070_gat), .Y(G2151_1122_gat) );
BUFX20 U_g1074 (.A(G1916_1077_gat), .Y(G1941_1123_gat) );
AND2XL U_g1075 (.A(G662_550_ngat), .B(G661_1080_ngat), .Y(G663_1124_gat) );
AND2XL U_g1076 (.A(G683_434_gat), .B(G681_1081_gat), .Y(G689_1125_gat) );
AND2XL U_g1077 (.A(G1656_552_gat), .B(G673_1082_gat), .Y(G1661_1126_gat) );
AND2XL U_g1078 (.A(G1609_577_gat), .B(G1539_1079_gat), .Y(G1612_1127_gat) );
AND2XL U_g1079 (.A(G1618_578_gat), .B(G1584_1083_gat), .Y(G1621_1128_gat) );
AND2XL U_g1080 (.A(G1627_579_gat), .B(G1588_1084_gat), .Y(G1630_1129_gat) );
AND2XL U_g1081 (.A(G1636_580_gat), .B(G1592_1085_gat), .Y(G1639_1130_gat) );
AND2XL U_g1082 (.A(G1645_581_gat), .B(G1596_1086_gat), .Y(G1648_1131_gat) );
AND2XL U_g1083 (.A(G1654_582_gat), .B(G1600_1087_gat), .Y(G1657_1132_gat) );
AND2XL U_g1084 (.A(G1663_583_gat), .B(G1604_1088_gat), .Y(G1666_1133_gat) );
AND2XL U_g1085 (.A(G1672_584_gat), .B(G1608_1089_gat), .Y(G1675_1134_gat) );
AND2XL U_g1086 (.A(G620_1093_gat), .B(G619_1091_gat), .Y(G356_1135_gat) );
AND2XL U_g1087 (.A(G583_1094_gat), .B(G582_1092_gat), .Y(G357_1136_gat) );
BUFX20 U_g1088 (.A(G2458_1096_gat), .Y(G2461_1137_gat) );
BUFX20 U_g1089 (.A(G2458_1096_gat), .Y(G3323_1138_gat) );
BUFX20 U_g1090 (.A(G2375_1097_gat), .Y(G3208_1139_gat) );
BUFX20 U_g1091 (.A(G2375_1097_gat), .Y(G3216_1140_gat) );
BUFX20 U_g1092 (.A(G2445_1098_gat), .Y(G2530_1141_gat) );
BUFX20 U_g1093 (.A(G2448_1099_gat), .Y(G2451_1142_gat) );
BUFX20 U_g1094 (.A(G2328_1101_gat), .Y(G3142_1143_gat) );
BUFX20 U_g1095 (.A(G2328_1101_gat), .Y(G3150_1144_gat) );
AND3XL U_g1096 (.A(G2151_1122_ngat), .B(G2150_1102_ngat), .C(G2149_1104_ngat), .Y(G2156_1145_gat) );
AND3XL U_g1097 (.A(G1941_1123_ngat), .B(G1940_1103_ngat), .C(G1939_1105_ngat), .Y(G1946_1146_gat) );
BUFX20 U_g1098 (.A(G2262_1106_gat), .Y(G2388_1147_gat) );
BUFX20 U_g1099 (.A(G2210_1107_gat), .Y(G2380_1148_gat) );
AND2XL U_g1100 (.A(G2146_1108_ngat), .B(G2143_1116_ngat), .Y(G2152_1149_gat) );
AND2XL U_g1101 (.A(G2146_1108_ngat), .B(G2143_1116_ngat), .Y(G2155_1150_gat) );
BUFX20 U_g1102 (.A(G2103_1110_gat), .Y(G2364_1151_gat) );
BUFX20 U_g1103 (.A(G2048_1111_gat), .Y(G2351_1152_gat) );
BUFX20 U_g1104 (.A(G1998_1112_gat), .Y(G2338_1153_gat) );
AND2XL U_g1105 (.A(G1936_1113_ngat), .B(G1933_1117_ngat), .Y(G1942_1154_gat) );
AND2XL U_g1106 (.A(G1936_1113_ngat), .B(G1933_1117_ngat), .Y(G1945_1155_gat) );
BUFX20 U_g1107 (.A(G1895_1115_gat), .Y(G2317_1156_gat) );
AND3XL U_g1108 (.A(G691_524_ngat), .B(G690_535_ngat), .C(G689_1125_ngat), .Y(G692_1157_gat) );
AND2XL U_g1109 (.A(G3070_1119_gat), .B(G3063_1013_gat), .Y(G607_1158_gat) );
AND2XL U_g1110 (.A(G3078_1121_gat), .B(G3071_1014_gat), .Y(G604_1159_gat) );
AND2XL U_g1111 (.A(G694_435_gat), .B(G663_1124_gat), .Y(G700_1160_gat) );
AND2XL U_g1112 (.A(G357_1136_gat), .B(G356_1135_gat), .Y(G358_1161_gat) );
BUFX20 U_g1113 (.A(G3323_1138_gat), .Y(G3329_1162_gat) );
BUFX20 U_g1114 (.A(G3208_1139_gat), .Y(G3212_1163_gat) );
BUFX20 U_g1115 (.A(G3216_1140_gat), .Y(G3220_1164_gat) );
AND2XL U_g1116 (.A(G2293_238_gat), .B(G2152_1149_gat), .Y(G2454_1165_gat) );
AND2XL U_g1117 (.A(G2288_240_gat), .B(G1942_1154_gat), .Y(G2444_1166_gat) );
BUFX20 U_g1118 (.A(G3142_1143_gat), .Y(G3146_1167_gat) );
BUFX20 U_g1119 (.A(G3150_1144_gat), .Y(G3154_1168_gat) );
AND2XL U_g1120 (.A(G2156_1145_gat), .B(G2155_1150_gat), .Y(G2157_1169_gat) );
AND2XL U_g1121 (.A(G1946_1146_gat), .B(G1945_1155_gat), .Y(G1947_1170_gat) );
BUFX20 U_g1122 (.A(G2388_1147_gat), .Y(G3237_1171_gat) );
BUFX20 U_g1123 (.A(G2388_1147_gat), .Y(G3245_1172_gat) );
BUFX20 U_g1124 (.A(G2380_1148_gat), .Y(G3221_1173_gat) );
BUFX20 U_g1125 (.A(G2380_1148_gat), .Y(G3229_1174_gat) );
AND2XL U_g1126 (.A(G2152_1149_gat), .B(G2103_1110_gat), .Y(G2312_1175_gat) );
BUFX20 U_g1127 (.A(G2364_1151_gat), .Y(G3187_1176_gat) );
BUFX20 U_g1128 (.A(G2364_1151_gat), .Y(G3197_1177_gat) );
BUFX20 U_g1129 (.A(G2351_1152_gat), .Y(G3171_1178_gat) );
BUFX20 U_g1130 (.A(G2351_1152_gat), .Y(G3179_1179_gat) );
BUFX20 U_g1131 (.A(G2338_1153_gat), .Y(G3155_1180_gat) );
BUFX20 U_g1132 (.A(G2338_1153_gat), .Y(G3163_1181_gat) );
AND2XL U_g1133 (.A(G1942_1154_gat), .B(G1895_1115_gat), .Y(G2272_1182_gat) );
BUFX20 U_g1134 (.A(G2317_1156_gat), .Y(G3121_1183_gat) );
BUFX20 U_g1135 (.A(G2317_1156_gat), .Y(G3131_1184_gat) );
AND2XL U_g1136 (.A(G607_1158_gat), .B(G606_1118_gat), .Y(G608_1185_gat) );
AND2XL U_g1137 (.A(G604_1159_gat), .B(G603_1120_gat), .Y(G605_1186_gat) );
AND3XL U_g1138 (.A(G702_530_ngat), .B(G701_523_ngat), .C(G700_1160_ngat), .Y(G703_1187_gat) );
AND2XL U_g1139 (.A(G1674_554_gat), .B(G692_1157_gat), .Y(G1679_1188_gat) );
AND2XL U_g1140 (.A(G3228_1040_gat), .B(G3221_1173_gat), .Y(G2432_1189_gat) );
AND2XL U_g1141 (.A(G3236_1041_gat), .B(G3229_1174_gat), .Y(G2387_1190_gat) );
AND2XL U_g1142 (.A(G3244_1042_gat), .B(G3237_1171_gat), .Y(G2395_1191_gat) );
AND2XL U_g1143 (.A(G3252_1043_gat), .B(G3245_1172_gat), .Y(G2400_1192_gat) );
BUFX20 U_g1144 (.A(G2454_1165_gat), .Y(G2533_1193_gat) );
AND2XL U_g1145 (.A(G3162_1044_gat), .B(G3155_1180_gat), .Y(G2345_1194_gat) );
AND2XL U_g1146 (.A(G3170_1045_gat), .B(G3163_1181_gat), .Y(G2350_1195_gat) );
AND2XL U_g1147 (.A(G3178_1046_gat), .B(G3171_1178_gat), .Y(G2358_1196_gat) );
AND2XL U_g1148 (.A(G3186_1047_gat), .B(G3179_1179_gat), .Y(G2363_1197_gat) );
AND2XL U_g1149 (.A(G3194_1048_gat), .B(G3187_1176_gat), .Y(G3196_1198_gat) );
AND2XL U_g1150 (.A(G3204_1049_gat), .B(G3197_1177_gat), .Y(G2371_1199_gat) );
BUFX20 U_g1151 (.A(G2444_1166_gat), .Y(G2523_1200_gat) );
AND2XL U_g1152 (.A(G3128_1050_gat), .B(G3121_1183_gat), .Y(G3130_1201_gat) );
AND2XL U_g1153 (.A(G3138_1051_gat), .B(G3131_1184_gat), .Y(G2324_1202_gat) );
BUFX20 U_g1154 (.A(G2157_1169_gat), .Y(G2372_1203_gat) );
BUFX20 U_g1155 (.A(G1947_1170_gat), .Y(G2325_1204_gat) );
AND4XL U_g1156 (.A(G2103_1110_gat), .B(G2210_1107_gat), .C(G2157_1169_gat), .D(G2257_1053_gat), .Y(G2314_1205_gat) );
AND4XL U_g1157 (.A(G2262_1106_gat), .B(G2210_1107_gat), .C(G2157_1169_gat), .D(G2103_1110_gat), .Y(G2309_1206_gat) );
BUFX20 U_g1158 (.A(G3237_1171_gat), .Y(G3243_1207_gat) );
BUFX20 U_g1159 (.A(G3245_1172_gat), .Y(G3251_1208_gat) );
AND3XL U_g1160 (.A(G2205_1055_gat), .B(G2157_1169_gat), .C(G2103_1110_gat), .Y(G2313_1209_gat) );
BUFX20 U_g1161 (.A(G3221_1173_gat), .Y(G3227_1210_gat) );
BUFX20 U_g1162 (.A(G3229_1174_gat), .Y(G3235_1211_gat) );
BUFX20 U_g1163 (.A(G3187_1176_gat), .Y(G3193_1212_gat) );
BUFX20 U_g1164 (.A(G3197_1177_gat), .Y(G3203_1213_gat) );
AND4XL U_g1165 (.A(G1895_1115_gat), .B(G1998_1112_gat), .C(G1947_1170_gat), .D(G2043_1059_gat), .Y(G2274_1214_gat) );
AND4XL U_g1166 (.A(G2048_1111_gat), .B(G1998_1112_gat), .C(G1947_1170_gat), .D(G1895_1115_gat), .Y(G2265_1215_gat) );
BUFX20 U_g1167 (.A(G3171_1178_gat), .Y(G3177_1216_gat) );
BUFX20 U_g1168 (.A(G3179_1179_gat), .Y(G3185_1217_gat) );
AND3XL U_g1169 (.A(G1993_1061_gat), .B(G1947_1170_gat), .C(G1895_1115_gat), .Y(G2273_1218_gat) );
BUFX20 U_g1170 (.A(G3155_1180_gat), .Y(G3161_1219_gat) );
BUFX20 U_g1171 (.A(G3163_1181_gat), .Y(G3169_1220_gat) );
BUFX20 U_g1172 (.A(G3121_1183_gat), .Y(G3127_1221_gat) );
BUFX20 U_g1173 (.A(G3131_1184_gat), .Y(G3137_1222_gat) );
BUFX20 U_g1174 (.A(G608_1185_gat), .Y(G350_1223_gat) );
BUFX20 U_g1175 (.A(G605_1186_gat), .Y(G349_1224_gat) );
AND2XL U_g1176 (.A(G1665_553_gat), .B(G703_1187_gat), .Y(G1670_1225_gat) );
AND2XL U_g1177 (.A(G3227_1210_gat), .B(G3224_975_gat), .Y(G2431_1226_gat) );
AND2XL U_g1178 (.A(G3235_1211_gat), .B(G3232_976_gat), .Y(G2386_1227_gat) );
AND2XL U_g1179 (.A(G3243_1207_gat), .B(G3240_977_gat), .Y(G2394_1228_gat) );
AND2XL U_g1180 (.A(G3251_1208_gat), .B(G3248_978_gat), .Y(G2399_1229_gat) );
AND2XL U_g1181 (.A(G2485_369_gat), .B(G2309_1206_gat), .Y(G2490_1230_gat) );
AND2XL U_g1182 (.A(G3161_1219_gat), .B(G3158_979_gat), .Y(G2344_1231_gat) );
AND2XL U_g1183 (.A(G3169_1220_gat), .B(G3166_980_gat), .Y(G2349_1232_gat) );
AND2XL U_g1184 (.A(G3177_1216_gat), .B(G3174_981_gat), .Y(G2357_1233_gat) );
AND2XL U_g1185 (.A(G3185_1217_gat), .B(G3182_982_gat), .Y(G2362_1234_gat) );
AND2XL U_g1186 (.A(G3193_1212_gat), .B(G3190_983_gat), .Y(G3195_1235_gat) );
AND2XL U_g1187 (.A(G3203_1213_gat), .B(G3200_984_gat), .Y(G2370_1236_gat) );
AND2XL U_g1188 (.A(G3127_1221_gat), .B(G3124_985_gat), .Y(G3129_1237_gat) );
AND2XL U_g1189 (.A(G3137_1222_gat), .B(G3134_986_gat), .Y(G2323_1238_gat) );
BUFX20 U_g1190 (.A(G2372_1203_gat), .Y(G3205_1239_gat) );
BUFX20 U_g1191 (.A(G2372_1203_gat), .Y(G3213_1240_gat) );
BUFX20 U_g1192 (.A(G2325_1204_gat), .Y(G3139_1241_gat) );
BUFX20 U_g1193 (.A(G2325_1204_gat), .Y(G3147_1242_gat) );
AND2XL U_g1194 (.A(G2265_1215_gat), .B(G2309_1206_gat), .Y(G372_1243_gat) );
AND4XL U_g1195 (.A(G2314_1205_gat), .B(G2313_1209_gat), .C(G2312_1175_gat), .D(G2311_1109_gat), .Y(G2315_1244_gat) );
BUFX20 U_g1196 (.A(G2265_1215_gat), .Y(G2268_1245_gat) );
AND4XL U_g1197 (.A(G2274_1214_gat), .B(G2273_1218_gat), .C(G2272_1182_gat), .D(G2271_1114_gat), .Y(G2275_1246_gat) );
AND2XL U_g1198 (.A(G350_1223_gat), .B(G349_1224_gat), .Y(G351_1247_gat) );
AND2XL U_g1199 (.A(G2302_236_gat), .B(G2315_1244_gat), .Y(G2464_1248_gat) );
AND2XL U_g1200 (.A(G3212_1163_gat), .B(G3205_1239_gat), .Y(G2425_1249_gat) );
AND2XL U_g1201 (.A(G3220_1164_gat), .B(G3213_1240_gat), .Y(G2379_1250_gat) );
AND2XL U_g1202 (.A(G2432_1189_gat), .B(G2431_1226_gat), .Y(G2433_1251_gat) );
AND2XL U_g1203 (.A(G2387_1190_gat), .B(G2386_1227_gat), .Y(G1669_1252_gat) );
AND2XL U_g1204 (.A(G2395_1191_gat), .B(G2394_1228_gat), .Y(G2396_1253_gat) );
AND2XL U_g1205 (.A(G2400_1192_gat), .B(G2399_1229_gat), .Y(G1678_1254_gat) );
AND2XL U_g1206 (.A(G2490_1230_ngat), .B(G2489_1100_ngat), .Y(G2491_1255_gat) );
AND2XL U_g1207 (.A(G2345_1194_gat), .B(G2344_1231_gat), .Y(G2346_1256_gat) );
AND2XL U_g1208 (.A(G2350_1195_gat), .B(G2349_1232_gat), .Y(G1633_1257_gat) );
AND2XL U_g1209 (.A(G2358_1196_gat), .B(G2357_1233_gat), .Y(G2359_1258_gat) );
AND2XL U_g1210 (.A(G2363_1197_gat), .B(G2362_1234_gat), .Y(G1642_1259_gat) );
AND2XL U_g1211 (.A(G3196_1198_gat), .B(G3195_1235_gat), .Y(G3308_1260_gat) );
AND2XL U_g1212 (.A(G2371_1199_gat), .B(G2370_1236_gat), .Y(G1651_1261_gat) );
AND2XL U_g1213 (.A(G3130_1201_gat), .B(G3129_1237_gat), .Y(G3272_1262_gat) );
AND2XL U_g1214 (.A(G2324_1202_gat), .B(G2323_1238_gat), .Y(G1615_1263_gat) );
AND2XL U_g1215 (.A(G3146_1167_gat), .B(G3139_1241_gat), .Y(G2332_1264_gat) );
AND2XL U_g1216 (.A(G3154_1168_gat), .B(G3147_1242_gat), .Y(G2337_1265_gat) );
BUFX20 U_g1217 (.A(G3205_1239_gat), .Y(G3211_1266_gat) );
BUFX20 U_g1218 (.A(G3213_1240_gat), .Y(G3219_1267_gat) );
BUFX20 U_g1219 (.A(G3139_1241_gat), .Y(G3145_1268_gat) );
BUFX20 U_g1220 (.A(G3147_1242_gat), .Y(G3153_1269_gat) );
AND2XL U_g1221 (.A(G2315_1244_gat), .B(G2265_1215_gat), .Y(G2307_1270_gat) );
BUFX20 U_g1222 (.A(G2275_1246_gat), .Y(G2308_1271_gat) );
AND2XL U_g1223 (.A(G2396_1253_gat), .B(G330_46_gat), .Y(G2612_1272_gat) );
AND2XL U_g1224 (.A(G2491_1255_gat), .B(G330_46_gat), .Y(G3374_1273_gat) );
AND2XL U_g1225 (.A(G2461_1137_gat), .B(G2433_1251_gat), .Y(G2518_1274_gat) );
BUFX20 U_g1226 (.A(G2464_1248_gat), .Y(G2467_1275_gat) );
BUFX20 U_g1227 (.A(G2464_1248_gat), .Y(G3295_1276_gat) );
AND2XL U_g1228 (.A(G3211_1266_gat), .B(G3208_1139_gat), .Y(G2424_1277_gat) );
AND2XL U_g1229 (.A(G3219_1267_gat), .B(G3216_1140_gat), .Y(G2378_1278_gat) );
BUFX20 U_g1230 (.A(G2433_1251_gat), .Y(G3326_1279_gat) );
BUFX20 U_g1231 (.A(G1669_1252_gat), .Y(G1667_1280_gat) );
BUFX20 U_g1232 (.A(G2396_1253_gat), .Y(G2439_1281_gat) );
BUFX20 U_g1233 (.A(G1678_1254_gat), .Y(G1676_1282_gat) );
BUFX20 U_g1234 (.A(G2491_1255_gat), .Y(G2495_1283_gat) );
BUFX20 U_g1235 (.A(G2346_1256_gat), .Y(G2406_1284_gat) );
BUFX20 U_g1236 (.A(G2346_1256_gat), .Y(G2409_1285_gat) );
BUFX20 U_g1237 (.A(G1633_1257_gat), .Y(G1631_1286_gat) );
BUFX20 U_g1238 (.A(G2359_1258_gat), .Y(G2415_1287_gat) );
BUFX20 U_g1239 (.A(G2359_1258_gat), .Y(G2419_1288_gat) );
BUFX20 U_g1240 (.A(G1642_1259_gat), .Y(G1640_1289_gat) );
BUFX20 U_g1241 (.A(G3308_1260_gat), .Y(G3312_1290_gat) );
BUFX20 U_g1242 (.A(G1651_1261_gat), .Y(G1649_1291_gat) );
BUFX20 U_g1243 (.A(G3272_1262_gat), .Y(G3276_1292_gat) );
BUFX20 U_g1244 (.A(G1615_1263_gat), .Y(G1613_1293_gat) );
AND2XL U_g1245 (.A(G3145_1268_gat), .B(G3142_1143_gat), .Y(G2331_1294_gat) );
AND2XL U_g1246 (.A(G3153_1269_gat), .B(G3150_1144_gat), .Y(G2336_1295_gat) );
AND2XL U_g1247 (.A(G2308_1271_gat), .B(G2307_1270_gat), .Y(G368_1296_gat) );
BUFX20 U_g1248 (.A(G2612_1272_gat), .Y(G3406_1297_gat) );
BUFX20 U_g1249 (.A(G2612_1272_gat), .Y(G3414_1298_gat) );
BUFX20 U_g1250 (.A(G3374_1273_gat), .Y(G3378_1299_gat) );
AND2XL U_g1251 (.A(G2518_1274_ngat), .B(G2455_1095_ngat), .Y(G2519_1300_gat) );
AND2XL U_g1252 (.A(G3329_1162_gat), .B(G3326_1279_gat), .Y(G2607_1301_gat) );
AND2XL U_g1253 (.A(G2415_1287_gat), .B(G2467_1275_gat), .Y(G2517_1302_gat) );
AND3XL U_g1254 (.A(G2467_1275_gat), .B(G2419_1288_gat), .C(G2409_1285_gat), .Y(G2532_1303_gat) );
BUFX20 U_g1255 (.A(G2467_1275_gat), .Y(G2642_1304_gat) );
BUFX20 U_g1256 (.A(G2467_1275_gat), .Y(G2645_1305_gat) );
BUFX20 U_g1257 (.A(G3295_1276_gat), .Y(G3301_1306_gat) );
AND2XL U_g1258 (.A(G2425_1249_gat), .B(G2424_1277_gat), .Y(G2426_1307_gat) );
AND2XL U_g1259 (.A(G2379_1250_gat), .B(G2378_1278_gat), .Y(G1660_1308_gat) );
AND2XL U_g1260 (.A(G2433_1251_gat), .B(G2439_1281_gat), .Y(G2514_1309_gat) );
BUFX20 U_g1261 (.A(G3326_1279_gat), .Y(G3330_1310_gat) );
AND2XL U_g1262 (.A(G2439_1281_gat), .B(G2439_1281_gat), .Y(G3422_1311_gat) );
AND2XL U_g1263 (.A(G2451_1142_gat), .B(G2409_1285_gat), .Y(G2531_1312_gat) );
AND3XL U_g1264 (.A(G2409_1285_gat), .B(G2419_1288_gat), .C(G2495_1283_gat), .Y(G2511_1313_gat) );
AND2XL U_g1265 (.A(G2415_1287_gat), .B(G2495_1283_gat), .Y(G2512_1314_gat) );
BUFX20 U_g1266 (.A(G2409_1285_gat), .Y(G3290_1315_gat) );
BUFX20 U_g1267 (.A(G2415_1287_gat), .Y(G3298_1316_gat) );
AND2XL U_g1268 (.A(G2332_1264_gat), .B(G2331_1294_gat), .Y(G2333_1317_gat) );
AND2XL U_g1269 (.A(G2337_1265_gat), .B(G2336_1295_gat), .Y(G1624_1318_gat) );
AND2XL U_g1270 (.A(G2268_1245_gat), .B(G2467_1275_gat), .Y(G2500_1319_gat) );
AND2XL U_g1271 (.A(G2268_1245_gat), .B(G2495_1283_gat), .Y(G2505_1320_gat) );
BUFX20 U_g1272 (.A(G368_1296_gat), .Y(G369_1321_gat) );
AND2XL U_g1273 (.A(G1646_436_gat), .B(G1649_1291_gat), .Y(G1650_1322_gat) );
AND2XL U_g1274 (.A(G1664_438_gat), .B(G1667_1280_gat), .Y(G1668_1323_gat) );
AND2XL U_g1275 (.A(G1673_439_gat), .B(G1676_1282_gat), .Y(G1677_1324_gat) );
AND2XL U_g1276 (.A(G1610_446_gat), .B(G1613_1293_gat), .Y(G1614_1325_gat) );
AND2XL U_g1277 (.A(G1628_448_gat), .B(G1631_1286_gat), .Y(G1632_1326_gat) );
AND2XL U_g1278 (.A(G1637_449_gat), .B(G1640_1289_gat), .Y(G1641_1327_gat) );
AND3XL U_g1279 (.A(G2642_1304_gat), .B(G2491_1255_gat), .C(G330_46_gat), .Y(G2643_1328_gat) );
AND2XL U_g1280 (.A(G3425_130_gat), .B(G3422_1311_gat), .Y(G2624_1329_gat) );
BUFX20 U_g1281 (.A(G3406_1297_gat), .Y(G3410_1330_gat) );
BUFX20 U_g1282 (.A(G3414_1298_gat), .Y(G3418_1331_gat) );
AND2XL U_g1283 (.A(G2514_1309_gat), .B(G330_46_gat), .Y(G3398_1332_gat) );
AND2XL U_g1284 (.A(G2512_1314_gat), .B(G330_46_gat), .Y(G2567_1333_gat) );
AND2XL U_g1285 (.A(G2511_1313_gat), .B(G330_46_gat), .Y(G3350_1334_gat) );
AND2XL U_g1286 (.A(G2455_1095_gat), .B(G2426_1307_gat), .Y(G2534_1335_gat) );
BUFX20 U_g1287 (.A(G2519_1300_gat), .Y(G3313_1336_gat) );
BUFX20 U_g1288 (.A(G2519_1300_gat), .Y(G2654_1337_gat) );
AND3XL U_g1289 (.A(G2461_1137_gat), .B(G2433_1251_gat), .C(G2426_1307_gat), .Y(G2535_1338_gat) );
AND2XL U_g1290 (.A(G3330_1310_gat), .B(G3323_1138_gat), .Y(G2608_1339_gat) );
AND2XL U_g1291 (.A(G3301_1306_gat), .B(G3298_1316_gat), .Y(G3303_1340_gat) );
BUFX20 U_g1292 (.A(G2426_1307_gat), .Y(G3316_1341_gat) );
BUFX20 U_g1293 (.A(G1660_1308_gat), .Y(G1658_1342_gat) );
AND3XL U_g1294 (.A(G2426_1307_gat), .B(G2433_1251_gat), .C(G2439_1281_gat), .Y(G2513_1343_gat) );
BUFX20 U_g1295 (.A(G3422_1311_gat), .Y(G3426_1344_gat) );
AND3XL U_g1296 (.A(G2532_1303_gat), .B(G2531_1312_gat), .C(G2530_1141_gat), .Y(G3277_1345_gat) );
AND2XL U_g1297 (.A(G2517_1302_ngat), .B(G2448_1099_ngat), .Y(G3287_1346_gat) );
BUFX20 U_g1298 (.A(G3290_1315_gat), .Y(G3294_1347_gat) );
BUFX20 U_g1299 (.A(G3298_1316_gat), .Y(G3302_1348_gat) );
BUFX20 U_g1300 (.A(G2333_1317_gat), .Y(G3280_1349_gat) );
BUFX20 U_g1301 (.A(G2333_1317_gat), .Y(G2401_1350_gat) );
BUFX20 U_g1302 (.A(G1624_1318_gat), .Y(G1622_1351_gat) );
BUFX20 U_g1303 (.A(G2505_1320_gat), .Y(G3253_1352_gat) );
AND2XL U_g1304 (.A(G2500_1319_ngat), .B(G2275_1246_ngat), .Y(G2501_1353_gat) );
AND3XL U_g1305 (.A(G1643_727_ngat), .B(G1641_1327_ngat), .C(G1639_1130_ngat), .Y(G1644_1354_gat) );
AND3XL U_g1306 (.A(G1634_730_ngat), .B(G1632_1326_ngat), .C(G1630_1129_ngat), .Y(G1635_1355_gat) );
AND3XL U_g1307 (.A(G1616_733_ngat), .B(G1614_1325_ngat), .C(G1612_1127_ngat), .Y(G1617_1356_gat) );
AND3XL U_g1308 (.A(G1652_1090_ngat), .B(G1650_1322_ngat), .C(G1648_1131_ngat), .Y(G1653_1357_gat) );
AND3XL U_g1309 (.A(G1670_1225_ngat), .B(G1668_1323_ngat), .C(G1666_1133_ngat), .Y(G1671_1358_gat) );
AND3XL U_g1310 (.A(G1679_1188_ngat), .B(G1677_1324_ngat), .C(G1675_1134_ngat), .Y(G1680_1359_gat) );
AND2XL U_g1311 (.A(G3426_1344_gat), .B(G3419_51_gat), .Y(G2625_1360_gat) );
BUFX20 U_g1312 (.A(G3398_1332_gat), .Y(G3402_1361_gat) );
AND2XL U_g1313 (.A(G2513_1343_gat), .B(G330_46_gat), .Y(G2589_1362_gat) );
BUFX20 U_g1314 (.A(G2567_1333_gat), .Y(G3358_1363_gat) );
BUFX20 U_g1315 (.A(G2567_1333_gat), .Y(G3366_1364_gat) );
BUFX20 U_g1316 (.A(G3350_1334_gat), .Y(G3354_1365_gat) );
AND2XL U_g1317 (.A(G2654_1337_gat), .B(G2519_1300_gat), .Y(G398_1366_gat) );
BUFX20 U_g1318 (.A(G3313_1336_gat), .Y(G3319_1367_gat) );
BUFX20 U_g1319 (.A(G2654_1337_gat), .Y(G2657_1368_gat) );
AND2XL U_g1320 (.A(G2608_1339_gat), .B(G2607_1301_gat), .Y(G2609_1369_gat) );
AND4XL U_g1321 (.A(G2467_1275_gat), .B(G2419_1288_gat), .C(G2406_1284_gat), .D(G2401_1350_gat), .Y(G2526_1370_gat) );
AND2XL U_g1322 (.A(G2645_1305_ngat), .B(G2643_1328_ngat), .Y(G932_1371_gat) );
AND2XL U_g1323 (.A(G2645_1305_ngat), .B(G2643_1328_ngat), .Y(G2647_1372_gat) );
AND2XL U_g1324 (.A(G3302_1348_gat), .B(G3295_1276_gat), .Y(G3304_1373_gat) );
BUFX20 U_g1325 (.A(G3316_1341_gat), .Y(G3320_1374_gat) );
AND2XL U_g1326 (.A(G2445_1098_gat), .B(G2401_1350_gat), .Y(G2524_1375_gat) );
BUFX20 U_g1327 (.A(G3277_1345_gat), .Y(G3283_1376_gat) );
AND3XL U_g1328 (.A(G2451_1142_gat), .B(G2406_1284_gat), .C(G2401_1350_gat), .Y(G2525_1377_gat) );
AND2XL U_g1329 (.A(G3294_1347_gat), .B(G3287_1346_gat), .Y(G2563_1378_gat) );
BUFX20 U_g1330 (.A(G3287_1346_gat), .Y(G3293_1379_gat) );
AND3XL U_g1331 (.A(G2535_1338_gat), .B(G2534_1335_gat), .C(G2533_1193_gat), .Y(G3305_1380_gat) );
AND4XL U_g1332 (.A(G2419_1288_gat), .B(G2409_1285_gat), .C(G2401_1350_gat), .D(G2495_1283_gat), .Y(G2508_1381_gat) );
BUFX20 U_g1333 (.A(G3280_1349_gat), .Y(G3284_1382_gat) );
BUFX20 U_g1334 (.A(G3253_1352_gat), .Y(G3259_1383_gat) );
BUFX20 U_g1335 (.A(G2501_1353_gat), .Y(G3264_1384_gat) );
BUFX20 U_g1336 (.A(G2501_1353_gat), .Y(G2629_1385_gat) );
AND2XL U_g1337 (.A(G1655_437_gat), .B(G1658_1342_gat), .Y(G1659_1386_gat) );
AND2XL U_g1338 (.A(G1619_447_gat), .B(G1622_1351_gat), .Y(G1623_1387_gat) );
AND2XL U_g1339 (.A(G2680_568_gat), .B(G1617_1356_gat), .Y(G2687_1388_gat) );
AND2XL U_g1340 (.A(G2718_570_gat), .B(G1635_1355_gat), .Y(G2725_1389_gat) );
AND2XL U_g1341 (.A(G2735_571_gat), .B(G1644_1354_gat), .Y(G2742_1390_gat) );
AND2XL U_g1342 (.A(G2753_572_gat), .B(G1653_1357_gat), .Y(G2760_1391_gat) );
AND2XL U_g1343 (.A(G2787_574_gat), .B(G1671_1358_gat), .Y(G2794_1392_gat) );
AND2XL U_g1344 (.A(G2804_575_gat), .B(G1680_1359_gat), .Y(G2811_1393_gat) );
AND3XL U_g1345 (.A(G2657_1368_gat), .B(G2514_1309_gat), .C(G330_46_gat), .Y(G397_1394_gat) );
AND2XL U_g1346 (.A(G2625_1360_gat), .B(G2624_1329_gat), .Y(G2626_1395_gat) );
BUFX20 U_g1347 (.A(G2589_1362_gat), .Y(G3382_1396_gat) );
BUFX20 U_g1348 (.A(G2589_1362_gat), .Y(G3390_1397_gat) );
BUFX20 U_g1349 (.A(G3358_1363_gat), .Y(G3362_1398_gat) );
BUFX20 U_g1350 (.A(G3366_1364_gat), .Y(G3370_1399_gat) );
AND2XL U_g1351 (.A(G2508_1381_gat), .B(G330_46_gat), .Y(G2544_1400_gat) );
AND2XL U_g1352 (.A(G3320_1374_gat), .B(G3313_1336_gat), .Y(G3322_1401_gat) );
BUFX20 U_g1353 (.A(G2609_1369_gat), .Y(G3403_1402_gat) );
BUFX20 U_g1354 (.A(G2609_1369_gat), .Y(G3411_1403_gat) );
BUFX20 U_g1355 (.A(G2647_1372_gat), .Y(G2650_1404_gat) );
AND2XL U_g1356 (.A(G3304_1373_gat), .B(G3303_1340_gat), .Y(G3371_1405_gat) );
AND2XL U_g1357 (.A(G3319_1367_gat), .B(G3316_1341_gat), .Y(G3321_1406_gat) );
AND2XL U_g1358 (.A(G3284_1382_gat), .B(G3277_1345_gat), .Y(G3286_1407_gat) );
BUFX20 U_g1359 (.A(G3305_1380_gat), .Y(G3311_1408_gat) );
BUFX20 U_g1360 (.A(G2508_1381_gat), .Y(G3256_1409_gat) );
AND2XL U_g1361 (.A(G3293_1379_gat), .B(G3290_1315_gat), .Y(G2562_1410_gat) );
AND2XL U_g1362 (.A(G3312_1290_gat), .B(G3305_1380_gat), .Y(G2585_1411_gat) );
AND4XL U_g1363 (.A(G2526_1370_gat), .B(G2525_1377_gat), .C(G2524_1375_gat), .D(G2523_1200_gat), .Y(G2527_1412_gat) );
AND2XL U_g1364 (.A(G3283_1376_gat), .B(G3280_1349_gat), .Y(G3285_1413_gat) );
BUFX20 U_g1365 (.A(G3264_1384_gat), .Y(G3268_1414_gat) );
BUFX20 U_g1366 (.A(G2629_1385_gat), .Y(G2632_1415_gat) );
AND2XL U_g1367 (.A(G2629_1385_gat), .B(G2501_1353_gat), .Y(G2634_1416_gat) );
AND3XL U_g1368 (.A(G1625_732_ngat), .B(G1623_1387_ngat), .C(G1621_1128_ngat), .Y(G1626_1417_gat) );
AND3XL U_g1369 (.A(G1661_1126_ngat), .B(G1659_1386_ngat), .C(G1657_1132_ngat), .Y(G1662_1418_gat) );
AND2XL U_g1370 (.A(G927_347_gat), .B(G932_1371_gat), .Y(G933_1419_gat) );
AND3XL U_g1371 (.A(G2632_1415_gat), .B(G2505_1320_gat), .C(G330_46_gat), .Y(G2633_1420_gat) );
AND2XL U_g1372 (.A(G3410_1330_gat), .B(G3403_1402_gat), .Y(G2616_1421_gat) );
AND2XL U_g1373 (.A(G3418_1331_gat), .B(G3411_1403_gat), .Y(G2622_1422_gat) );
BUFX20 U_g1374 (.A(G3382_1396_gat), .Y(G3386_1423_gat) );
BUFX20 U_g1375 (.A(G3390_1397_gat), .Y(G3394_1424_gat) );
AND2XL U_g1376 (.A(G3378_1299_gat), .B(G3371_1405_gat), .Y(G2580_1425_gat) );
BUFX20 U_g1377 (.A(G2544_1400_gat), .Y(G3334_1426_gat) );
BUFX20 U_g1378 (.A(G2544_1400_gat), .Y(G3342_1427_gat) );
AND2XL U_g1379 (.A(G398_1366_ngat), .B(G397_1394_ngat), .Y(G399_1428_gat) );
AND2XL U_g1380 (.A(G3322_1401_gat), .B(G3321_1406_gat), .Y(G3395_1429_gat) );
BUFX20 U_g1381 (.A(G3403_1402_gat), .Y(G3409_1430_gat) );
BUFX20 U_g1382 (.A(G3411_1403_gat), .Y(G3417_1431_gat) );
BUFX20 U_g1383 (.A(G2650_1404_gat), .Y(G3454_1432_gat) );
BUFX20 U_g1384 (.A(G3371_1405_gat), .Y(G3377_1433_gat) );
AND2XL U_g1385 (.A(G3286_1407_gat), .B(G3285_1413_gat), .Y(G3347_1434_gat) );
AND2XL U_g1386 (.A(G2563_1378_gat), .B(G2562_1410_gat), .Y(G2564_1435_gat) );
BUFX20 U_g1387 (.A(G3256_1409_gat), .Y(G3260_1436_gat) );
AND2XL U_g1388 (.A(G3311_1408_gat), .B(G3308_1260_gat), .Y(G2584_1437_gat) );
BUFX20 U_g1389 (.A(G2527_1412_gat), .Y(G3261_1438_gat) );
BUFX20 U_g1390 (.A(G2527_1412_gat), .Y(G3269_1439_gat) );
AND2XL U_g1391 (.A(G3259_1383_gat), .B(G3256_1409_gat), .Y(G2536_1440_gat) );
AND3XL U_g1392 (.A(G938_722_ngat), .B(G933_1419_ngat), .C(G929_734_ngat), .Y(G362_1441_gat) );
AND3XL U_g1393 (.A(G938_722_ngat), .B(G933_1419_ngat), .C(G929_734_ngat), .Y(G1030_1442_gat) );
AND2XL U_g1394 (.A(G2803_562_gat), .B(G2626_1395_gat), .Y(G2808_1443_gat) );
AND2XL U_g1395 (.A(G2699_569_gat), .B(G1626_1417_gat), .Y(G2706_1444_gat) );
AND2XL U_g1396 (.A(G2770_573_gat), .B(G1662_1418_gat), .Y(G2777_1445_gat) );
AND2XL U_g1397 (.A(G2802_469_gat), .B(G2626_1395_gat), .Y(G2805_1446_gat) );
AND2XL U_g1398 (.A(G3409_1430_gat), .B(G3406_1297_gat), .Y(G2615_1447_gat) );
AND2XL U_g1399 (.A(G3417_1431_gat), .B(G3414_1298_gat), .Y(G2621_1448_gat) );
AND2XL U_g1400 (.A(G3402_1361_gat), .B(G3395_1429_gat), .Y(G2602_1449_gat) );
AND2XL U_g1401 (.A(G3377_1433_gat), .B(G3374_1273_gat), .Y(G2579_1450_gat) );
AND2XL U_g1402 (.A(G3354_1365_gat), .B(G3347_1434_gat), .Y(G2557_1451_gat) );
BUFX20 U_g1403 (.A(G3334_1426_gat), .Y(G3338_1452_gat) );
BUFX20 U_g1404 (.A(G3342_1427_gat), .Y(G3346_1453_gat) );
BUFX20 U_g1405 (.A(G3395_1429_gat), .Y(G3401_1454_gat) );
BUFX20 U_g1406 (.A(G3454_1432_gat), .Y(G3458_1455_gat) );
BUFX20 U_g1407 (.A(G3347_1434_gat), .Y(G3353_1456_gat) );
BUFX20 U_g1408 (.A(G2564_1435_gat), .Y(G3355_1457_gat) );
BUFX20 U_g1409 (.A(G2564_1435_gat), .Y(G3363_1458_gat) );
AND2XL U_g1410 (.A(G2585_1411_gat), .B(G2584_1437_gat), .Y(G2586_1459_gat) );
BUFX20 U_g1411 (.A(G3261_1438_gat), .Y(G3267_1460_gat) );
BUFX20 U_g1412 (.A(G3269_1439_gat), .Y(G3275_1461_gat) );
AND2XL U_g1413 (.A(G3276_1292_gat), .B(G3269_1439_gat), .Y(G2540_1462_gat) );
AND2XL U_g1414 (.A(G3260_1436_gat), .B(G3253_1352_gat), .Y(G2537_1463_gat) );
AND2XL U_g1415 (.A(G3268_1414_gat), .B(G3261_1438_gat), .Y(G3112_1464_gat) );
AND2XL U_g1416 (.A(G2634_1416_ngat), .B(G2633_1420_ngat), .Y(G2635_1465_gat) );
BUFX20 U_g1417 (.A(G1030_1442_gat), .Y(G363_1466_gat) );
AND3XL U_g1418 (.A(G2811_1393_ngat), .B(G2808_1443_ngat), .C(G2805_1446_ngat), .Y(G2814_1467_gat) );
AND3XL U_g1419 (.A(G2811_1393_ngat), .B(G2808_1443_ngat), .C(G2805_1446_ngat), .Y(G2816_1468_gat) );
AND2XL U_g1420 (.A(G2616_1421_gat), .B(G2615_1447_gat), .Y(G2617_1469_gat) );
AND2XL U_g1421 (.A(G2622_1422_gat), .B(G2621_1448_gat), .Y(G2623_1470_gat) );
AND2XL U_g1422 (.A(G3401_1454_gat), .B(G3398_1332_gat), .Y(G2601_1471_gat) );
AND2XL U_g1423 (.A(G2580_1425_gat), .B(G2579_1450_gat), .Y(G2581_1472_gat) );
AND2XL U_g1424 (.A(G3362_1398_gat), .B(G3355_1457_gat), .Y(G2571_1473_gat) );
AND2XL U_g1425 (.A(G3370_1399_gat), .B(G3363_1458_gat), .Y(G2577_1474_gat) );
AND2XL U_g1426 (.A(G3353_1456_gat), .B(G3350_1334_gat), .Y(G2556_1475_gat) );
BUFX20 U_g1427 (.A(G3355_1457_gat), .Y(G3361_1476_gat) );
BUFX20 U_g1428 (.A(G3363_1458_gat), .Y(G3369_1477_gat) );
BUFX20 U_g1429 (.A(G2586_1459_gat), .Y(G3379_1478_gat) );
BUFX20 U_g1430 (.A(G2586_1459_gat), .Y(G3387_1479_gat) );
AND2XL U_g1431 (.A(G3275_1461_gat), .B(G3272_1262_gat), .Y(G2539_1480_gat) );
AND2XL U_g1432 (.A(G2537_1463_gat), .B(G2536_1440_gat), .Y(G2538_1481_gat) );
AND2XL U_g1433 (.A(G3267_1460_gat), .B(G3264_1384_gat), .Y(G3111_1482_gat) );
BUFX20 U_g1434 (.A(G2635_1465_gat), .Y(G2638_1483_gat) );
AND2XL U_g1435 (.A(G363_1466_gat), .B(G362_1441_gat), .Y(G364_1484_gat) );
BUFX20 U_g1436 (.A(G2814_1467_gat), .Y(G3459_1485_gat) );
BUFX20 U_g1437 (.A(G2816_1468_gat), .Y(G395_1486_gat) );
BUFX20 U_g1438 (.A(G2623_1470_gat), .Y(G3451_1487_gat) );
AND2XL U_g1439 (.A(G2602_1449_gat), .B(G2601_1471_gat), .Y(G2603_1488_gat) );
AND2XL U_g1440 (.A(G3386_1423_gat), .B(G3379_1478_gat), .Y(G2593_1489_gat) );
AND2XL U_g1441 (.A(G3394_1424_gat), .B(G3387_1479_gat), .Y(G2598_1490_gat) );
AND2XL U_g1442 (.A(G3361_1476_gat), .B(G3358_1363_gat), .Y(G2570_1491_gat) );
AND2XL U_g1443 (.A(G3369_1477_gat), .B(G3366_1364_gat), .Y(G2576_1492_gat) );
AND2XL U_g1444 (.A(G2557_1451_gat), .B(G2556_1475_gat), .Y(G2558_1493_gat) );
AND2XL U_g1445 (.A(G2538_1481_gat), .B(G330_46_gat), .Y(G3116_1494_gat) );
AND2XL U_g1446 (.A(G2647_1372_gat), .B(G2617_1469_gat), .Y(G3446_1495_gat) );
BUFX20 U_g1447 (.A(G3379_1478_gat), .Y(G3385_1496_gat) );
BUFX20 U_g1448 (.A(G3387_1479_gat), .Y(G3393_1497_gat) );
AND2XL U_g1449 (.A(G2540_1462_gat), .B(G2539_1480_gat), .Y(G2541_1498_gat) );
AND2XL U_g1450 (.A(G3112_1464_gat), .B(G3111_1482_gat), .Y(G3113_1499_gat) );
BUFX20 U_g1451 (.A(G2638_1483_gat), .Y(G3438_1500_gat) );
AND2XL U_g1452 (.A(G2734_558_gat), .B(G2581_1472_gat), .Y(G2739_1501_gat) );
AND2XL U_g1453 (.A(G2733_465_gat), .B(G2581_1472_gat), .Y(G2736_1502_gat) );
AND2XL U_g1454 (.A(G2785_468_gat), .B(G2617_1469_gat), .Y(G2788_1503_gat) );
AND2XL U_g1455 (.A(G395_1486_gat), .B(G2814_1467_gat), .Y(G396_1504_gat) );
BUFX20 U_g1456 (.A(G3459_1485_gat), .Y(G3465_1505_gat) );
BUFX20 U_g1457 (.A(G3451_1487_gat), .Y(G3457_1506_gat) );
BUFX20 U_g1458 (.A(G2603_1488_gat), .Y(G3443_1507_gat) );
AND2XL U_g1459 (.A(G3385_1496_gat), .B(G3382_1396_gat), .Y(G2592_1508_gat) );
AND2XL U_g1460 (.A(G3393_1497_gat), .B(G3390_1397_gat), .Y(G2597_1509_gat) );
AND2XL U_g1461 (.A(G2571_1473_gat), .B(G2570_1491_gat), .Y(G2572_1510_gat) );
AND2XL U_g1462 (.A(G2577_1474_gat), .B(G2576_1492_gat), .Y(G2578_1511_gat) );
BUFX20 U_g1463 (.A(G2558_1493_gat), .Y(G3427_1512_gat) );
BUFX20 U_g1464 (.A(G3116_1494_gat), .Y(G3120_1513_gat) );
AND2XL U_g1465 (.A(G3458_1455_gat), .B(G3451_1487_gat), .Y(G2677_1514_gat) );
BUFX20 U_g1466 (.A(G3446_1495_gat), .Y(G3450_1515_gat) );
BUFX20 U_g1467 (.A(G2541_1498_gat), .Y(G3331_1516_gat) );
BUFX20 U_g1468 (.A(G2541_1498_gat), .Y(G3339_1517_gat) );
BUFX20 U_g1469 (.A(G3113_1499_gat), .Y(G3119_1518_gat) );
BUFX20 U_g1470 (.A(G3438_1500_gat), .Y(G3442_1519_gat) );
AND2XL U_g1471 (.A(G2697_463_gat), .B(G2558_1493_gat), .Y(G2700_1520_gat) );
AND3XL U_g1472 (.A(G2742_1390_ngat), .B(G2739_1501_ngat), .C(G2736_1502_ngat), .Y(G2745_1521_gat) );
AND3XL U_g1473 (.A(G2742_1390_ngat), .B(G2739_1501_ngat), .C(G2736_1502_ngat), .Y(G2748_1522_gat) );
AND2XL U_g1474 (.A(G2768_467_gat), .B(G2603_1488_gat), .Y(G2771_1523_gat) );
AND2XL U_g1475 (.A(G3450_1515_gat), .B(G3443_1507_gat), .Y(G2672_1524_gat) );
BUFX20 U_g1476 (.A(G3443_1507_gat), .Y(G3449_1525_gat) );
AND2XL U_g1477 (.A(G2593_1489_gat), .B(G2592_1508_gat), .Y(G2594_1526_gat) );
AND2XL U_g1478 (.A(G2598_1490_gat), .B(G2597_1509_gat), .Y(G2599_1527_gat) );
BUFX20 U_g1479 (.A(G2578_1511_gat), .Y(G3435_1528_gat) );
BUFX20 U_g1480 (.A(G3427_1512_gat), .Y(G3433_1529_gat) );
AND2XL U_g1481 (.A(G3338_1452_gat), .B(G3331_1516_gat), .Y(G2548_1530_gat) );
AND2XL U_g1482 (.A(G3346_1453_gat), .B(G3339_1517_gat), .Y(G2553_1531_gat) );
AND2XL U_g1483 (.A(G3119_1518_gat), .B(G3116_1494_gat), .Y(G954_1532_gat) );
AND2XL U_g1484 (.A(G3457_1506_gat), .B(G3454_1432_gat), .Y(G2676_1533_gat) );
BUFX20 U_g1485 (.A(G3331_1516_gat), .Y(G3337_1534_gat) );
BUFX20 U_g1486 (.A(G3339_1517_gat), .Y(G3345_1535_gat) );
AND2XL U_g1487 (.A(G3120_1513_gat), .B(G3113_1499_gat), .Y(G955_1536_gat) );
AND2XL U_g1488 (.A(G2635_1465_gat), .B(G2572_1510_gat), .Y(G3430_1537_gat) );
AND2XL U_g1489 (.A(G2716_464_gat), .B(G2572_1510_gat), .Y(G2719_1538_gat) );
BUFX20 U_g1490 (.A(G2745_1521_gat), .Y(G3491_1539_gat) );
BUFX20 U_g1491 (.A(G2745_1521_gat), .Y(G3499_1540_gat) );
BUFX20 U_g1492 (.A(G2748_1522_gat), .Y(G383_1541_gat) );
BUFX20 U_g1493 (.A(G2599_1527_gat), .Y(G2600_1542_gat) );
BUFX20 U_g1494 (.A(G3435_1528_gat), .Y(G3441_1543_gat) );
AND2XL U_g1495 (.A(G3433_1529_gat), .B(G3430_1537_gat), .Y(G2664_1544_gat) );
AND2XL U_g1496 (.A(G3337_1534_gat), .B(G3334_1426_gat), .Y(G2547_1545_gat) );
AND2XL U_g1497 (.A(G3345_1535_gat), .B(G3342_1427_gat), .Y(G2552_1546_gat) );
AND2XL U_g1498 (.A(G955_1536_gat), .B(G954_1532_gat), .Y(G950_1547_gat) );
AND4XL U_g1499 (.A(G2650_1404_gat), .B(G2594_1526_gat), .C(G2603_1488_gat), .D(G2617_1469_gat), .Y(G2662_1548_gat) );
AND2XL U_g1500 (.A(G2677_1514_gat), .B(G2676_1533_gat), .Y(G2674_1549_gat) );
AND2XL U_g1501 (.A(G3449_1525_gat), .B(G3446_1495_gat), .Y(G2671_1550_gat) );
AND2XL U_g1502 (.A(G3442_1519_gat), .B(G3435_1528_gat), .Y(G2670_1551_gat) );
BUFX20 U_g1503 (.A(G3430_1537_gat), .Y(G3434_1552_gat) );
AND2XL U_g1504 (.A(G383_1541_gat), .B(G2745_1521_gat), .Y(G384_1553_gat) );
BUFX20 U_g1505 (.A(G3491_1539_gat), .Y(G3497_1554_gat) );
BUFX20 U_g1506 (.A(G3499_1540_gat), .Y(G3505_1555_gat) );
AND2XL U_g1507 (.A(G2751_466_gat), .B(G2594_1526_gat), .Y(G2754_1556_gat) );
AND2XL U_g1508 (.A(G2672_1524_gat), .B(G2671_1550_gat), .Y(G2673_1557_gat) );
AND2XL U_g1509 (.A(G3434_1552_gat), .B(G3427_1512_gat), .Y(G2665_1558_gat) );
AND2XL U_g1510 (.A(G2548_1530_gat), .B(G2547_1545_gat), .Y(G2549_1559_gat) );
AND2XL U_g1511 (.A(G2553_1531_gat), .B(G2552_1546_gat), .Y(G2554_1560_gat) );
AND2XL U_g1512 (.A(G2650_1404_ngat), .B(G2600_1542_ngat), .Y(G2661_1561_gat) );
BUFX20 U_g1513 (.A(G2674_1549_gat), .Y(G2675_1562_gat) );
AND2XL U_g1514 (.A(G3441_1543_gat), .B(G3438_1500_gat), .Y(G2669_1563_gat) );
AND2XL U_g1515 (.A(G943_445_gat), .B(G950_1547_gat), .Y(G951_1564_gat) );
AND2XL U_g1516 (.A(G2665_1558_gat), .B(G2664_1544_gat), .Y(G2666_1565_gat) );
BUFX20 U_g1517 (.A(G2554_1560_gat), .Y(G2555_1566_gat) );
AND2XL U_g1518 (.A(G2662_1548_ngat), .B(G2661_1561_ngat), .Y(G2663_1567_gat) );
AND4XL U_g1519 (.A(G2638_1483_gat), .B(G2549_1559_gat), .C(G2558_1493_gat), .D(G2572_1510_gat), .Y(G2659_1568_gat) );
AND2XL U_g1520 (.A(G2670_1551_gat), .B(G2669_1563_gat), .Y(G2667_1569_gat) );
AND3XL U_g1521 (.A(G951_1564_ngat), .B(G947_910_ngat), .C(G944_969_ngat), .Y(G365_1570_gat) );
AND3XL U_g1522 (.A(G951_1564_ngat), .B(G947_910_ngat), .C(G944_969_ngat), .Y(G1031_1571_gat) );
AND2XL U_g1523 (.A(G2769_560_gat), .B(G2673_1557_gat), .Y(G2774_1572_gat) );
AND2XL U_g1524 (.A(G2786_561_gat), .B(G2675_1562_gat), .Y(G2791_1573_gat) );
AND2XL U_g1525 (.A(G2678_462_gat), .B(G2549_1559_gat), .Y(G2681_1574_gat) );
AND2XL U_g1526 (.A(G2638_1483_ngat), .B(G2555_1566_ngat), .Y(G2658_1575_gat) );
BUFX20 U_g1527 (.A(G2667_1569_gat), .Y(G2668_1576_gat) );
BUFX20 U_g1528 (.A(G1031_1571_gat), .Y(G366_1577_gat) );
AND2XL U_g1529 (.A(G2698_556_gat), .B(G2666_1565_gat), .Y(G2703_1578_gat) );
AND2XL U_g1530 (.A(G2752_559_gat), .B(G2663_1567_gat), .Y(G2757_1579_gat) );
AND3XL U_g1531 (.A(G2777_1445_ngat), .B(G2774_1572_ngat), .C(G2771_1523_ngat), .Y(G2780_1580_gat) );
AND3XL U_g1532 (.A(G2777_1445_ngat), .B(G2774_1572_ngat), .C(G2771_1523_ngat), .Y(G2782_1581_gat) );
AND3XL U_g1533 (.A(G2794_1392_ngat), .B(G2791_1573_ngat), .C(G2788_1503_ngat), .Y(G2797_1582_gat) );
AND3XL U_g1534 (.A(G2794_1392_ngat), .B(G2791_1573_ngat), .C(G2788_1503_ngat), .Y(G2799_1583_gat) );
AND2XL U_g1535 (.A(G2659_1568_ngat), .B(G2658_1575_ngat), .Y(G2660_1584_gat) );
AND2XL U_g1536 (.A(G366_1577_gat), .B(G365_1570_gat), .Y(G367_1585_gat) );
AND2XL U_g1537 (.A(G2717_557_gat), .B(G2668_1576_gat), .Y(G2722_1586_gat) );
AND3XL U_g1538 (.A(G2706_1444_ngat), .B(G2703_1578_ngat), .C(G2700_1520_ngat), .Y(G2709_1587_gat) );
AND3XL U_g1539 (.A(G2706_1444_ngat), .B(G2703_1578_ngat), .C(G2700_1520_ngat), .Y(G2713_1588_gat) );
AND3XL U_g1540 (.A(G2760_1391_ngat), .B(G2757_1579_ngat), .C(G2754_1556_ngat), .Y(G2763_1589_gat) );
AND3XL U_g1541 (.A(G2760_1391_ngat), .B(G2757_1579_ngat), .C(G2754_1556_ngat), .Y(G2765_1590_gat) );
BUFX20 U_g1542 (.A(G2780_1580_gat), .Y(G3467_1591_gat) );
BUFX20 U_g1543 (.A(G2782_1581_gat), .Y(G389_1592_gat) );
BUFX20 U_g1544 (.A(G2797_1582_gat), .Y(G3462_1593_gat) );
BUFX20 U_g1545 (.A(G2799_1583_gat), .Y(G392_1594_gat) );
AND2XL U_g1546 (.A(G2871_128_gat), .B(G2709_1587_gat), .Y(G2883_1595_gat) );
AND2XL U_g1547 (.A(G2679_555_gat), .B(G2660_1584_gat), .Y(G2684_1596_gat) );
AND2XL U_g1548 (.A(G2709_1587_gat), .B(G2709_1587_gat), .Y(G378_1597_gat) );
BUFX20 U_g1549 (.A(G2709_1587_gat), .Y(G3507_1598_gat) );
AND3XL U_g1550 (.A(G2725_1389_ngat), .B(G2722_1586_ngat), .C(G2719_1538_ngat), .Y(G2728_1599_gat) );
AND3XL U_g1551 (.A(G2725_1389_ngat), .B(G2722_1586_ngat), .C(G2719_1538_ngat), .Y(G2730_1600_gat) );
BUFX20 U_g1552 (.A(G2763_1589_gat), .Y(G3470_1601_gat) );
BUFX20 U_g1553 (.A(G2765_1590_gat), .Y(G386_1602_gat) );
AND2XL U_g1554 (.A(G389_1592_gat), .B(G2780_1580_gat), .Y(G390_1603_gat) );
BUFX20 U_g1555 (.A(G3467_1591_gat), .Y(G3473_1604_gat) );
AND2XL U_g1556 (.A(G392_1594_gat), .B(G2797_1582_gat), .Y(G393_1605_gat) );
BUFX20 U_g1557 (.A(G3462_1593_gat), .Y(G3466_1606_gat) );
AND2XL U_g1558 (.A(G3465_1505_gat), .B(G3462_1593_gat), .Y(G2821_1607_gat) );
AND4XL U_g1559 (.A(G2765_1590_gat), .B(G2782_1581_gat), .C(G2799_1583_gat), .D(G2816_1468_gat), .Y(G2922_1608_gat) );
BUFX20 U_g1560 (.A(G2883_1595_gat), .Y(G3544_1609_gat) );
BUFX20 U_g1561 (.A(G2883_1595_gat), .Y(G3552_1610_gat) );
AND3XL U_g1562 (.A(G2687_1388_ngat), .B(G2684_1596_ngat), .C(G2681_1574_ngat), .Y(G2690_1611_gat) );
AND3XL U_g1563 (.A(G2687_1388_ngat), .B(G2684_1596_ngat), .C(G2681_1574_ngat), .Y(G2694_1612_gat) );
BUFX20 U_g1564 (.A(G3507_1598_gat), .Y(G3513_1613_gat) );
BUFX20 U_g1565 (.A(G2728_1599_gat), .Y(G2839_1614_gat) );
BUFX20 U_g1566 (.A(G2730_1600_gat), .Y(G380_1615_gat) );
AND2XL U_g1567 (.A(G386_1602_gat), .B(G2763_1589_gat), .Y(G387_1616_gat) );
AND2XL U_g1568 (.A(G3473_1604_gat), .B(G3470_1601_gat), .Y(G2826_1617_gat) );
BUFX20 U_g1569 (.A(G3470_1601_gat), .Y(G3474_1618_gat) );
AND2XL U_g1570 (.A(G3466_1606_gat), .B(G3459_1485_gat), .Y(G2822_1619_gat) );
AND2XL U_g1571 (.A(G2690_1611_gat), .B(G2871_128_gat), .Y(G2880_1620_gat) );
BUFX20 U_g1572 (.A(G3544_1609_gat), .Y(G3548_1621_gat) );
BUFX20 U_g1573 (.A(G3552_1610_gat), .Y(G3556_1622_gat) );
AND3XL U_g1574 (.A(G2874_129_gat), .B(G2694_1612_gat), .C(G2713_1588_gat), .Y(G2928_1623_gat) );
AND2XL U_g1575 (.A(G2690_1611_gat), .B(G2690_1611_gat), .Y(G375_1624_gat) );
BUFX20 U_g1576 (.A(G2690_1611_gat), .Y(G3510_1625_gat) );
AND2XL U_g1577 (.A(G380_1615_gat), .B(G2728_1599_gat), .Y(G381_1626_gat) );
BUFX20 U_g1578 (.A(G2839_1614_gat), .Y(G3494_1627_gat) );
BUFX20 U_g1579 (.A(G2839_1614_gat), .Y(G3502_1628_gat) );
AND4XL U_g1580 (.A(G2694_1612_gat), .B(G2713_1588_gat), .C(G2730_1600_gat), .D(G2748_1522_gat), .Y(G2925_1629_gat) );
AND2XL U_g1581 (.A(G3474_1618_gat), .B(G3467_1591_gat), .Y(G2827_1630_gat) );
AND2XL U_g1582 (.A(G2822_1619_gat), .B(G2821_1607_gat), .Y(G2823_1631_gat) );
BUFX20 U_g1583 (.A(G2880_1620_gat), .Y(G3541_1632_gat) );
BUFX20 U_g1584 (.A(G2880_1620_gat), .Y(G3549_1633_gat) );
BUFX20 U_g1585 (.A(G3510_1625_gat), .Y(G3514_1634_gat) );
AND2XL U_g1586 (.A(G3513_1613_gat), .B(G3510_1625_gat), .Y(G3515_1635_gat) );
BUFX20 U_g1587 (.A(G3494_1627_gat), .Y(G3498_1636_gat) );
BUFX20 U_g1588 (.A(G3502_1628_gat), .Y(G3506_1637_gat) );
AND2XL U_g1589 (.A(G3497_1554_gat), .B(G3494_1627_gat), .Y(G2842_1638_gat) );
AND2XL U_g1590 (.A(G3505_1555_gat), .B(G3502_1628_gat), .Y(G2852_1639_gat) );
AND2XL U_g1591 (.A(G2827_1630_gat), .B(G2826_1617_gat), .Y(G2828_1640_gat) );
BUFX20 U_g1592 (.A(G2823_1631_gat), .Y(G3475_1641_gat) );
BUFX20 U_g1593 (.A(G2823_1631_gat), .Y(G3483_1642_gat) );
AND2XL U_g1594 (.A(G2925_1629_gat), .B(G2922_1608_gat), .Y(G406_1643_gat) );
AND2XL U_g1595 (.A(G2925_1629_gat), .B(G2922_1608_gat), .Y(G2929_1644_gat) );
BUFX20 U_g1596 (.A(G3541_1632_gat), .Y(G3547_1645_gat) );
BUFX20 U_g1597 (.A(G3549_1633_gat), .Y(G3555_1646_gat) );
AND2XL U_g1598 (.A(G3548_1621_gat), .B(G3541_1632_gat), .Y(G2887_1647_gat) );
AND2XL U_g1599 (.A(G3556_1622_gat), .B(G3549_1633_gat), .Y(G2896_1648_gat) );
AND2XL U_g1600 (.A(G2929_1644_ngat), .B(G2928_1623_ngat), .Y(G2930_1649_gat) );
AND2XL U_g1601 (.A(G3514_1634_gat), .B(G3507_1598_gat), .Y(G3516_1650_gat) );
AND2XL U_g1602 (.A(G3498_1636_gat), .B(G3491_1539_gat), .Y(G2843_1651_gat) );
AND2XL U_g1603 (.A(G3506_1637_gat), .B(G3499_1540_gat), .Y(G2853_1652_gat) );
BUFX20 U_g1604 (.A(G2828_1640_gat), .Y(G3478_1653_gat) );
BUFX20 U_g1605 (.A(G2828_1640_gat), .Y(G3486_1654_gat) );
BUFX20 U_g1606 (.A(G3475_1641_gat), .Y(G3481_1655_gat) );
BUFX20 U_g1607 (.A(G3483_1642_gat), .Y(G3489_1656_gat) );
BUFX20 U_g1608 (.A(G406_1643_gat), .Y(G407_1657_gat) );
AND2XL U_g1609 (.A(G3547_1645_gat), .B(G3544_1609_gat), .Y(G2886_1658_gat) );
AND2XL U_g1610 (.A(G3555_1646_gat), .B(G3552_1610_gat), .Y(G2895_1659_gat) );
AND2XL U_g1611 (.A(G2930_1649_gat), .B(G213_26_gat), .Y(G408_1660_gat) );
AND2XL U_g1612 (.A(G3516_1650_gat), .B(G3515_1635_gat), .Y(G3520_1661_gat) );
AND2XL U_g1613 (.A(G2843_1651_gat), .B(G2842_1638_gat), .Y(G2844_1662_gat) );
AND2XL U_g1614 (.A(G2853_1652_gat), .B(G2852_1639_gat), .Y(G2848_1663_gat) );
AND2XL U_g1615 (.A(G3481_1655_gat), .B(G3478_1653_gat), .Y(G2831_1664_gat) );
BUFX20 U_g1616 (.A(G3478_1653_gat), .Y(G3482_1665_gat) );
AND2XL U_g1617 (.A(G3489_1656_gat), .B(G3486_1654_gat), .Y(G2836_1666_gat) );
BUFX20 U_g1618 (.A(G3486_1654_gat), .Y(G3490_1667_gat) );
AND2XL U_g1619 (.A(G2887_1647_gat), .B(G2886_1658_gat), .Y(G2888_1668_gat) );
AND2XL U_g1620 (.A(G2896_1648_gat), .B(G2895_1659_gat), .Y(G2891_1669_gat) );
BUFX20 U_g1621 (.A(G408_1660_gat), .Y(G409_1670_gat) );
BUFX20 U_g1622 (.A(G3520_1661_gat), .Y(G3524_1671_gat) );
BUFX20 U_g1623 (.A(G2844_1662_gat), .Y(G3517_1672_gat) );
BUFX20 U_g1624 (.A(G2848_1663_gat), .Y(G2849_1673_gat) );
AND2XL U_g1625 (.A(G3482_1665_gat), .B(G3475_1641_gat), .Y(G2832_1674_gat) );
AND2XL U_g1626 (.A(G3490_1667_gat), .B(G3483_1642_gat), .Y(G2837_1675_gat) );
AND3XL U_g1627 (.A(G2903_349_gat), .B(G2888_1668_gat), .C(G2849_1673_gat), .Y(G2908_1676_gat) );
AND3XL U_g1628 (.A(G2900_350_gat), .B(G2888_1668_gat), .C(G2844_1662_gat), .Y(G2906_1677_gat) );
BUFX20 U_g1629 (.A(G2891_1669_gat), .Y(G2892_1678_gat) );
AND2XL U_g1630 (.A(G3524_1671_gat), .B(G3517_1672_gat), .Y(G2855_1679_gat) );
BUFX20 U_g1631 (.A(G3517_1672_gat), .Y(G3523_1680_gat) );
AND2XL U_g1632 (.A(G2832_1674_gat), .B(G2831_1664_gat), .Y(G2833_1681_gat) );
AND2XL U_g1633 (.A(G2837_1675_gat), .B(G2836_1666_gat), .Y(G2838_1682_gat) );
AND3XL U_g1634 (.A(G2903_349_gat), .B(G2892_1678_gat), .C(G2844_1662_gat), .Y(G2907_1683_gat) );
AND3XL U_g1635 (.A(G2900_350_gat), .B(G2892_1678_gat), .C(G2849_1673_gat), .Y(G2909_1684_gat) );
AND2XL U_g1636 (.A(G3523_1680_gat), .B(G3520_1661_gat), .Y(G2854_1685_gat) );
BUFX20 U_g1637 (.A(G2833_1681_gat), .Y(G3525_1686_gat) );
BUFX20 U_g1638 (.A(G2833_1681_gat), .Y(G3533_1687_gat) );
BUFX20 U_g1639 (.A(G2838_1682_gat), .Y(G2913_1688_gat) );
AND4XL U_g1640 (.A(G2909_1684_ngat), .B(G2908_1676_ngat), .C(G2907_1683_ngat), .D(G2906_1677_ngat), .Y(G2910_1689_gat) );
AND2XL U_g1641 (.A(G2855_1679_gat), .B(G2854_1685_gat), .Y(G2856_1690_gat) );
BUFX20 U_g1642 (.A(G3525_1686_gat), .Y(G3531_1691_gat) );
BUFX20 U_g1643 (.A(G3533_1687_gat), .Y(G3539_1692_gat) );
BUFX20 U_g1644 (.A(G2913_1688_gat), .Y(G3560_1693_gat) );
BUFX20 U_g1645 (.A(G2913_1688_gat), .Y(G3568_1694_gat) );
BUFX20 U_g1646 (.A(G2910_1689_gat), .Y(G3557_1695_gat) );
BUFX20 U_g1647 (.A(G2910_1689_gat), .Y(G3565_1696_gat) );
BUFX20 U_g1648 (.A(G2856_1690_gat), .Y(G3528_1697_gat) );
BUFX20 U_g1649 (.A(G2856_1690_gat), .Y(G3536_1698_gat) );
BUFX20 U_g1650 (.A(G3560_1693_gat), .Y(G3564_1699_gat) );
BUFX20 U_g1651 (.A(G3568_1694_gat), .Y(G3572_1700_gat) );
AND2XL U_g1652 (.A(G3564_1699_gat), .B(G3557_1695_gat), .Y(G2921_1701_gat) );
BUFX20 U_g1653 (.A(G3557_1695_gat), .Y(G3563_1702_gat) );
AND2XL U_g1654 (.A(G3572_1700_gat), .B(G3565_1696_gat), .Y(G2917_1703_gat) );
BUFX20 U_g1655 (.A(G3565_1696_gat), .Y(G3571_1704_gat) );
BUFX20 U_g1656 (.A(G3528_1697_gat), .Y(G3532_1705_gat) );
BUFX20 U_g1657 (.A(G3536_1698_gat), .Y(G3540_1706_gat) );
AND2XL U_g1658 (.A(G3531_1691_gat), .B(G3528_1697_gat), .Y(G2863_1707_gat) );
AND2XL U_g1659 (.A(G3539_1692_gat), .B(G3536_1698_gat), .Y(G2859_1708_gat) );
AND2XL U_g1660 (.A(G3532_1705_gat), .B(G3525_1686_gat), .Y(G2864_1709_gat) );
AND2XL U_g1661 (.A(G3540_1706_gat), .B(G3533_1687_gat), .Y(G2860_1710_gat) );
AND2XL U_g1662 (.A(G3563_1702_gat), .B(G3560_1693_gat), .Y(G2920_1711_gat) );
AND2XL U_g1663 (.A(G3571_1704_gat), .B(G3568_1694_gat), .Y(G2916_1712_gat) );
AND2XL U_g1664 (.A(G2921_1701_gat), .B(G2920_1711_gat), .Y(G403_1713_gat) );
AND2XL U_g1665 (.A(G2917_1703_gat), .B(G2916_1712_gat), .Y(G404_1714_gat) );
AND2XL U_g1666 (.A(G2864_1709_gat), .B(G2863_1707_gat), .Y(G400_1715_gat) );
AND2XL U_g1667 (.A(G2860_1710_gat), .B(G2859_1708_gat), .Y(G401_1716_gat) );
AND2XL U_g1668 (.A(G404_1714_gat), .B(G403_1713_gat), .Y(G405_1717_gat) );
AND2XL U_g1669 (.A(G401_1716_gat), .B(G400_1715_gat), .Y(G402_1718_gat) );
INVXL U_g1670 (.A(G257_34_gat), .Y(G257_34_ngat) );
INVXL U_g1671 (.A(G264_35_gat), .Y(G264_35_ngat) );
INVXL U_g1672 (.A(G41_4_gat), .Y(G41_4_ngat) );
INVXL U_g1673 (.A(G45_5_gat), .Y(G45_5_ngat) );
INVXL U_g1674 (.A(G1698_48_gat), .Y(G1698_48_ngat) );
INVXL U_g1675 (.A(G33_3_gat), .Y(G33_3_ngat) );
INVXL U_g1676 (.A(G2865_61_gat), .Y(G2865_61_ngat) );
INVXL U_g1677 (.A(G2868_50_gat), .Y(G2868_50_ngat) );
INVXL U_g1678 (.A(G1032_115_gat), .Y(G1032_115_ngat) );
INVXL U_g1679 (.A(G1035_63_gat), .Y(G1035_63_ngat) );
INVXL U_g1680 (.A(G1540_111_gat), .Y(G1540_111_ngat) );
INVXL U_g1681 (.A(G169_22_gat), .Y(G169_22_ngat) );
INVXL U_g1682 (.A(G758_108_gat), .Y(G758_108_ngat) );
INVXL U_g1683 (.A(G20_2_gat), .Y(G20_2_ngat) );
INVXL U_g1684 (.A(G2051_104_gat), .Y(G2051_104_ngat) );
INVXL U_g1685 (.A(G1_0_gat), .Y(G1_0_ngat) );
INVXL U_g1686 (.A(G1828_110_gat), .Y(G1828_110_ngat) );
INVXL U_g1687 (.A(G1772_212_gat), .Y(G1772_212_ngat) );
INVXL U_g1688 (.A(G116_13_gat), .Y(G116_13_ngat) );
INVXL U_g1689 (.A(G1773_345_gat), .Y(G1773_345_ngat) );
INVXL U_g1690 (.A(G107_12_gat), .Y(G107_12_ngat) );
INVXL U_g1691 (.A(G97_11_gat), .Y(G97_11_ngat) );
INVXL U_g1692 (.A(G87_10_gat), .Y(G87_10_ngat) );
INVXL U_g1693 (.A(G77_9_gat), .Y(G77_9_ngat) );
INVXL U_g1694 (.A(G68_8_gat), .Y(G68_8_ngat) );
INVXL U_g1695 (.A(G58_7_gat), .Y(G58_7_ngat) );
INVXL U_g1696 (.A(G50_6_gat), .Y(G50_6_ngat) );
INVXL U_g1697 (.A(G1768_351_gat), .Y(G1768_351_ngat) );
INVXL U_g1698 (.A(G1769_221_gat), .Y(G1769_221_ngat) );
INVXL U_g1699 (.A(G1770_357_gat), .Y(G1770_357_ngat) );
INVXL U_g1700 (.A(G1761_352_gat), .Y(G1761_352_ngat) );
INVXL U_g1701 (.A(G1762_223_gat), .Y(G1762_223_ngat) );
INVXL U_g1702 (.A(G1763_358_gat), .Y(G1763_358_ngat) );
INVXL U_g1703 (.A(G1754_353_gat), .Y(G1754_353_ngat) );
INVXL U_g1704 (.A(G1755_225_gat), .Y(G1755_225_ngat) );
INVXL U_g1705 (.A(G1756_360_gat), .Y(G1756_360_ngat) );
INVXL U_g1706 (.A(G1747_381_gat), .Y(G1747_381_ngat) );
INVXL U_g1707 (.A(G1748_228_gat), .Y(G1748_228_ngat) );
INVXL U_g1708 (.A(G1749_362_gat), .Y(G1749_362_ngat) );
INVXL U_g1709 (.A(G1740_385_gat), .Y(G1740_385_ngat) );
INVXL U_g1710 (.A(G1741_230_gat), .Y(G1741_230_ngat) );
INVXL U_g1711 (.A(G1742_364_gat), .Y(G1742_364_ngat) );
INVXL U_g1712 (.A(G1733_389_gat), .Y(G1733_389_ngat) );
INVXL U_g1713 (.A(G1734_232_gat), .Y(G1734_232_ngat) );
INVXL U_g1714 (.A(G1735_365_gat), .Y(G1735_365_ngat) );
INVXL U_g1715 (.A(G1726_396_gat), .Y(G1726_396_ngat) );
INVXL U_g1716 (.A(G1727_234_gat), .Y(G1727_234_ngat) );
INVXL U_g1717 (.A(G1728_367_gat), .Y(G1728_367_ngat) );
INVXL U_g1718 (.A(G1719_402_gat), .Y(G1719_402_ngat) );
INVXL U_g1719 (.A(G1720_235_gat), .Y(G1720_235_ngat) );
INVXL U_g1720 (.A(G1721_368_gat), .Y(G1721_368_ngat) );
INVXL U_g1721 (.A(G1025_244_gat), .Y(G1025_244_ngat) );
INVXL U_g1722 (.A(G1026_354_gat), .Y(G1026_354_ngat) );
INVXL U_g1723 (.A(G1027_393_gat), .Y(G1027_393_ngat) );
INVXL U_g1724 (.A(G1004_252_gat), .Y(G1004_252_ngat) );
INVXL U_g1725 (.A(G1005_392_gat), .Y(G1005_392_ngat) );
INVXL U_g1726 (.A(G1006_409_gat), .Y(G1006_409_ngat) );
INVXL U_g1727 (.A(G1018_253_gat), .Y(G1018_253_ngat) );
INVXL U_g1728 (.A(G1019_382_gat), .Y(G1019_382_ngat) );
INVXL U_g1729 (.A(G1020_398_gat), .Y(G1020_398_ngat) );
INVXL U_g1730 (.A(G997_259_gat), .Y(G997_259_ngat) );
INVXL U_g1731 (.A(G998_397_gat), .Y(G998_397_ngat) );
INVXL U_g1732 (.A(G999_415_gat), .Y(G999_415_ngat) );
INVXL U_g1733 (.A(G976_266_gat), .Y(G976_266_ngat) );
INVXL U_g1734 (.A(G977_414_gat), .Y(G977_414_ngat) );
INVXL U_g1735 (.A(G978_379_gat), .Y(G978_379_ngat) );
INVXL U_g1736 (.A(G990_267_gat), .Y(G990_267_ngat) );
INVXL U_g1737 (.A(G991_404_gat), .Y(G991_404_ngat) );
INVXL U_g1738 (.A(G992_418_gat), .Y(G992_418_ngat) );
INVXL U_g1739 (.A(G917_549_gat), .Y(G917_549_ngat) );
INVXL U_g1740 (.A(G920_361_gat), .Y(G920_361_ngat) );
INVXL U_g1741 (.A(G923_482_gat), .Y(G923_482_ngat) );
INVXL U_g1742 (.A(G2234_480_gat), .Y(G2234_480_ngat) );
INVXL U_g1743 (.A(G2235_472_gat), .Y(G2235_472_ngat) );
INVXL U_g1744 (.A(G2236_748_gat), .Y(G2236_748_ngat) );
INVXL U_g1745 (.A(G2182_483_gat), .Y(G2182_483_ngat) );
INVXL U_g1746 (.A(G2183_473_gat), .Y(G2183_473_ngat) );
INVXL U_g1747 (.A(G2184_747_gat), .Y(G2184_747_ngat) );
INVXL U_g1748 (.A(G2129_484_gat), .Y(G2129_484_ngat) );
INVXL U_g1749 (.A(G2130_474_gat), .Y(G2130_474_ngat) );
INVXL U_g1750 (.A(G2131_746_gat), .Y(G2131_746_ngat) );
INVXL U_g1751 (.A(G2077_487_gat), .Y(G2077_487_ngat) );
INVXL U_g1752 (.A(G2078_475_gat), .Y(G2078_475_ngat) );
INVXL U_g1753 (.A(G2079_745_gat), .Y(G2079_745_ngat) );
INVXL U_g1754 (.A(G2022_489_gat), .Y(G2022_489_ngat) );
INVXL U_g1755 (.A(G2023_476_gat), .Y(G2023_476_ngat) );
INVXL U_g1756 (.A(G2024_744_gat), .Y(G2024_744_ngat) );
INVXL U_g1757 (.A(G1972_493_gat), .Y(G1972_493_ngat) );
INVXL U_g1758 (.A(G1973_477_gat), .Y(G1973_477_ngat) );
INVXL U_g1759 (.A(G1974_743_gat), .Y(G1974_743_ngat) );
INVXL U_g1760 (.A(G1921_495_gat), .Y(G1921_495_ngat) );
INVXL U_g1761 (.A(G1922_478_gat), .Y(G1922_478_ngat) );
INVXL U_g1762 (.A(G1923_742_gat), .Y(G1923_742_ngat) );
INVXL U_g1763 (.A(G1871_499_gat), .Y(G1871_499_ngat) );
INVXL U_g1764 (.A(G1872_479_gat), .Y(G1872_479_ngat) );
INVXL U_g1765 (.A(G1873_741_gat), .Y(G1873_741_ngat) );
INVXL U_g1766 (.A(G2216_740_gat), .Y(G2216_740_ngat) );
INVXL U_g1767 (.A(G2219_380_gat), .Y(G2219_380_ngat) );
INVXL U_g1768 (.A(G2222_520_gat), .Y(G2222_520_ngat) );
INVXL U_g1769 (.A(G2164_739_gat), .Y(G2164_739_ngat) );
INVXL U_g1770 (.A(G2167_384_gat), .Y(G2167_384_ngat) );
INVXL U_g1771 (.A(G2170_525_gat), .Y(G2170_525_ngat) );
INVXL U_g1772 (.A(G2059_738_gat), .Y(G2059_738_ngat) );
INVXL U_g1773 (.A(G2062_395_gat), .Y(G2062_395_ngat) );
INVXL U_g1774 (.A(G2065_534_gat), .Y(G2065_534_ngat) );
INVXL U_g1775 (.A(G2004_737_gat), .Y(G2004_737_ngat) );
INVXL U_g1776 (.A(G2007_401_gat), .Y(G2007_401_ngat) );
INVXL U_g1777 (.A(G2010_537_gat), .Y(G2010_537_ngat) );
INVXL U_g1778 (.A(G1954_736_gat), .Y(G1954_736_ngat) );
INVXL U_g1779 (.A(G1957_407_gat), .Y(G1957_407_ngat) );
INVXL U_g1780 (.A(G1960_540_gat), .Y(G1960_540_ngat) );
INVXL U_g1781 (.A(G641_728_gat), .Y(G641_728_ngat) );
INVXL U_g1782 (.A(G644_269_gat), .Y(G644_269_ngat) );
INVXL U_g1783 (.A(G1853_735_gat), .Y(G1853_735_ngat) );
INVXL U_g1784 (.A(G1856_417_gat), .Y(G1856_417_ngat) );
INVXL U_g1785 (.A(G1859_547_gat), .Y(G1859_547_ngat) );
INVXL U_g1786 (.A(G1503_749_gat), .Y(G1503_749_ngat) );
INVXL U_g1787 (.A(G1504_777_gat), .Y(G1504_777_ngat) );
INVXL U_g1788 (.A(G1505_770_gat), .Y(G1505_770_ngat) );
INVXL U_g1789 (.A(G1506_764_gat), .Y(G1506_764_ngat) );
INVXL U_g1790 (.A(G1507_759_gat), .Y(G1507_759_ngat) );
INVXL U_g1791 (.A(G1508_755_gat), .Y(G1508_755_ngat) );
INVXL U_g1792 (.A(G1509_752_gat), .Y(G1509_752_ngat) );
INVXL U_g1793 (.A(G1510_750_gat), .Y(G1510_750_ngat) );
INVXL U_g1794 (.A(G1486_751_gat), .Y(G1486_751_ngat) );
INVXL U_g1795 (.A(G1487_844_gat), .Y(G1487_844_ngat) );
INVXL U_g1796 (.A(G1488_778_gat), .Y(G1488_778_ngat) );
INVXL U_g1797 (.A(G1489_771_gat), .Y(G1489_771_ngat) );
INVXL U_g1798 (.A(G1490_765_gat), .Y(G1490_765_ngat) );
INVXL U_g1799 (.A(G1491_760_gat), .Y(G1491_760_ngat) );
INVXL U_g1800 (.A(G1492_756_gat), .Y(G1492_756_ngat) );
INVXL U_g1801 (.A(G1493_753_gat), .Y(G1493_753_ngat) );
INVXL U_g1802 (.A(G1469_754_gat), .Y(G1469_754_ngat) );
INVXL U_g1803 (.A(G1470_853_gat), .Y(G1470_853_ngat) );
INVXL U_g1804 (.A(G1471_843_gat), .Y(G1471_843_ngat) );
INVXL U_g1805 (.A(G1472_779_gat), .Y(G1472_779_ngat) );
INVXL U_g1806 (.A(G1473_772_gat), .Y(G1473_772_ngat) );
INVXL U_g1807 (.A(G1474_766_gat), .Y(G1474_766_ngat) );
INVXL U_g1808 (.A(G1475_761_gat), .Y(G1475_761_ngat) );
INVXL U_g1809 (.A(G1476_757_gat), .Y(G1476_757_ngat) );
INVXL U_g1810 (.A(G1452_758_gat), .Y(G1452_758_ngat) );
INVXL U_g1811 (.A(G1453_861_gat), .Y(G1453_861_ngat) );
INVXL U_g1812 (.A(G1454_852_gat), .Y(G1454_852_ngat) );
INVXL U_g1813 (.A(G1455_842_gat), .Y(G1455_842_ngat) );
INVXL U_g1814 (.A(G1456_780_gat), .Y(G1456_780_ngat) );
INVXL U_g1815 (.A(G1457_773_gat), .Y(G1457_773_ngat) );
INVXL U_g1816 (.A(G1458_767_gat), .Y(G1458_767_ngat) );
INVXL U_g1817 (.A(G1459_762_gat), .Y(G1459_762_ngat) );
INVXL U_g1818 (.A(G1435_763_gat), .Y(G1435_763_ngat) );
INVXL U_g1819 (.A(G1436_870_gat), .Y(G1436_870_ngat) );
INVXL U_g1820 (.A(G1437_860_gat), .Y(G1437_860_ngat) );
INVXL U_g1821 (.A(G1438_851_gat), .Y(G1438_851_ngat) );
INVXL U_g1822 (.A(G1439_841_gat), .Y(G1439_841_ngat) );
INVXL U_g1823 (.A(G1440_781_gat), .Y(G1440_781_ngat) );
INVXL U_g1824 (.A(G1441_774_gat), .Y(G1441_774_ngat) );
INVXL U_g1825 (.A(G1442_768_gat), .Y(G1442_768_ngat) );
INVXL U_g1826 (.A(G1418_769_gat), .Y(G1418_769_ngat) );
INVXL U_g1827 (.A(G1419_879_gat), .Y(G1419_879_ngat) );
INVXL U_g1828 (.A(G1420_869_gat), .Y(G1420_869_ngat) );
INVXL U_g1829 (.A(G1421_859_gat), .Y(G1421_859_ngat) );
INVXL U_g1830 (.A(G1422_850_gat), .Y(G1422_850_ngat) );
INVXL U_g1831 (.A(G1423_840_gat), .Y(G1423_840_ngat) );
INVXL U_g1832 (.A(G1424_782_gat), .Y(G1424_782_ngat) );
INVXL U_g1833 (.A(G1425_775_gat), .Y(G1425_775_ngat) );
INVXL U_g1834 (.A(G1401_776_gat), .Y(G1401_776_ngat) );
INVXL U_g1835 (.A(G1402_889_gat), .Y(G1402_889_ngat) );
INVXL U_g1836 (.A(G1403_878_gat), .Y(G1403_878_ngat) );
INVXL U_g1837 (.A(G1404_868_gat), .Y(G1404_868_ngat) );
INVXL U_g1838 (.A(G1405_858_gat), .Y(G1405_858_ngat) );
INVXL U_g1839 (.A(G1406_849_gat), .Y(G1406_849_ngat) );
INVXL U_g1840 (.A(G1407_839_gat), .Y(G1407_839_ngat) );
INVXL U_g1841 (.A(G1408_783_gat), .Y(G1408_783_ngat) );
INVXL U_g1842 (.A(G1384_784_gat), .Y(G1384_784_ngat) );
INVXL U_g1843 (.A(G1385_898_gat), .Y(G1385_898_ngat) );
INVXL U_g1844 (.A(G1386_888_gat), .Y(G1386_888_ngat) );
INVXL U_g1845 (.A(G1387_877_gat), .Y(G1387_877_ngat) );
INVXL U_g1846 (.A(G1388_867_gat), .Y(G1388_867_ngat) );
INVXL U_g1847 (.A(G1389_857_gat), .Y(G1389_857_ngat) );
INVXL U_g1848 (.A(G1390_848_gat), .Y(G1390_848_ngat) );
INVXL U_g1849 (.A(G1391_838_gat), .Y(G1391_838_ngat) );
INVXL U_g1850 (.A(G1367_799_gat), .Y(G1367_799_ngat) );
INVXL U_g1851 (.A(G1368_847_gat), .Y(G1368_847_ngat) );
INVXL U_g1852 (.A(G1369_856_gat), .Y(G1369_856_ngat) );
INVXL U_g1853 (.A(G1370_866_gat), .Y(G1370_866_ngat) );
INVXL U_g1854 (.A(G1371_876_gat), .Y(G1371_876_ngat) );
INVXL U_g1855 (.A(G1372_887_gat), .Y(G1372_887_ngat) );
INVXL U_g1856 (.A(G1373_897_gat), .Y(G1373_897_ngat) );
INVXL U_g1857 (.A(G1374_907_gat), .Y(G1374_907_ngat) );
INVXL U_g1858 (.A(G1350_807_gat), .Y(G1350_807_ngat) );
INVXL U_g1859 (.A(G1351_855_gat), .Y(G1351_855_ngat) );
INVXL U_g1860 (.A(G1352_865_gat), .Y(G1352_865_ngat) );
INVXL U_g1861 (.A(G1353_875_gat), .Y(G1353_875_ngat) );
INVXL U_g1862 (.A(G1354_886_gat), .Y(G1354_886_ngat) );
INVXL U_g1863 (.A(G1355_896_gat), .Y(G1355_896_ngat) );
INVXL U_g1864 (.A(G1356_906_gat), .Y(G1356_906_ngat) );
INVXL U_g1865 (.A(G1357_800_gat), .Y(G1357_800_ngat) );
INVXL U_g1866 (.A(G1333_814_gat), .Y(G1333_814_ngat) );
INVXL U_g1867 (.A(G1334_864_gat), .Y(G1334_864_ngat) );
INVXL U_g1868 (.A(G1335_874_gat), .Y(G1335_874_ngat) );
INVXL U_g1869 (.A(G1336_885_gat), .Y(G1336_885_ngat) );
INVXL U_g1870 (.A(G1337_895_gat), .Y(G1337_895_ngat) );
INVXL U_g1871 (.A(G1338_905_gat), .Y(G1338_905_ngat) );
INVXL U_g1872 (.A(G1339_801_gat), .Y(G1339_801_ngat) );
INVXL U_g1873 (.A(G1340_808_gat), .Y(G1340_808_ngat) );
INVXL U_g1874 (.A(G1316_820_gat), .Y(G1316_820_ngat) );
INVXL U_g1875 (.A(G1317_873_gat), .Y(G1317_873_ngat) );
INVXL U_g1876 (.A(G1318_884_gat), .Y(G1318_884_ngat) );
INVXL U_g1877 (.A(G1319_894_gat), .Y(G1319_894_ngat) );
INVXL U_g1878 (.A(G1320_904_gat), .Y(G1320_904_ngat) );
INVXL U_g1879 (.A(G1321_802_gat), .Y(G1321_802_ngat) );
INVXL U_g1880 (.A(G1322_809_gat), .Y(G1322_809_ngat) );
INVXL U_g1881 (.A(G1323_815_gat), .Y(G1323_815_ngat) );
INVXL U_g1882 (.A(G1299_825_gat), .Y(G1299_825_ngat) );
INVXL U_g1883 (.A(G1300_883_gat), .Y(G1300_883_ngat) );
INVXL U_g1884 (.A(G1301_893_gat), .Y(G1301_893_ngat) );
INVXL U_g1885 (.A(G1302_903_gat), .Y(G1302_903_ngat) );
INVXL U_g1886 (.A(G1303_803_gat), .Y(G1303_803_ngat) );
INVXL U_g1887 (.A(G1304_810_gat), .Y(G1304_810_ngat) );
INVXL U_g1888 (.A(G1305_816_gat), .Y(G1305_816_ngat) );
INVXL U_g1889 (.A(G1306_821_gat), .Y(G1306_821_ngat) );
INVXL U_g1890 (.A(G1282_829_gat), .Y(G1282_829_ngat) );
INVXL U_g1891 (.A(G1283_892_gat), .Y(G1283_892_ngat) );
INVXL U_g1892 (.A(G1284_902_gat), .Y(G1284_902_ngat) );
INVXL U_g1893 (.A(G1285_804_gat), .Y(G1285_804_ngat) );
INVXL U_g1894 (.A(G1286_811_gat), .Y(G1286_811_ngat) );
INVXL U_g1895 (.A(G1287_817_gat), .Y(G1287_817_ngat) );
INVXL U_g1896 (.A(G1288_822_gat), .Y(G1288_822_ngat) );
INVXL U_g1897 (.A(G1289_826_gat), .Y(G1289_826_ngat) );
INVXL U_g1898 (.A(G1265_832_gat), .Y(G1265_832_ngat) );
INVXL U_g1899 (.A(G1266_901_gat), .Y(G1266_901_ngat) );
INVXL U_g1900 (.A(G1267_805_gat), .Y(G1267_805_ngat) );
INVXL U_g1901 (.A(G1268_812_gat), .Y(G1268_812_ngat) );
INVXL U_g1902 (.A(G1269_818_gat), .Y(G1269_818_ngat) );
INVXL U_g1903 (.A(G1270_823_gat), .Y(G1270_823_ngat) );
INVXL U_g1904 (.A(G1271_827_gat), .Y(G1271_827_ngat) );
INVXL U_g1905 (.A(G1272_830_gat), .Y(G1272_830_ngat) );
INVXL U_g1906 (.A(G1248_834_gat), .Y(G1248_834_ngat) );
INVXL U_g1907 (.A(G1249_806_gat), .Y(G1249_806_ngat) );
INVXL U_g1908 (.A(G1250_813_gat), .Y(G1250_813_ngat) );
INVXL U_g1909 (.A(G1251_819_gat), .Y(G1251_819_ngat) );
INVXL U_g1910 (.A(G1252_824_gat), .Y(G1252_824_ngat) );
INVXL U_g1911 (.A(G1253_828_gat), .Y(G1253_828_ngat) );
INVXL U_g1912 (.A(G1254_831_gat), .Y(G1254_831_ngat) );
INVXL U_g1913 (.A(G1255_833_gat), .Y(G1255_833_ngat) );
INVXL U_g1914 (.A(G983_908_gat), .Y(G983_908_ngat) );
INVXL U_g1915 (.A(G984_408_gat), .Y(G984_408_ngat) );
INVXL U_g1916 (.A(G985_378_gat), .Y(G985_378_ngat) );
INVXL U_g1917 (.A(G1011_909_gat), .Y(G1011_909_ngat) );
INVXL U_g1918 (.A(G1012_386_gat), .Y(G1012_386_ngat) );
INVXL U_g1919 (.A(G1013_403_gat), .Y(G1013_403_ngat) );
INVXL U_g1920 (.A(G614_968_gat), .Y(G614_968_ngat) );
INVXL U_g1921 (.A(G616_424_gat), .Y(G616_424_ngat) );
INVXL U_g1922 (.A(G617_536_gat), .Y(G617_536_ngat) );
INVXL U_g1923 (.A(G2482_949_gat), .Y(G2482_949_ngat) );
INVXL U_g1924 (.A(G2483_999_gat), .Y(G2483_999_ngat) );
INVXL U_g1925 (.A(G2248_1006_gat), .Y(G2248_1006_ngat) );
INVXL U_g1926 (.A(G2251_1000_gat), .Y(G2251_1000_ngat) );
INVXL U_g1927 (.A(G2196_1007_gat), .Y(G2196_1007_ngat) );
INVXL U_g1928 (.A(G2199_1001_gat), .Y(G2199_1001_ngat) );
INVXL U_g1929 (.A(G2091_1008_gat), .Y(G2091_1008_ngat) );
INVXL U_g1930 (.A(G2094_1002_gat), .Y(G2094_1002_ngat) );
INVXL U_g1931 (.A(G2034_1009_gat), .Y(G2034_1009_ngat) );
INVXL U_g1932 (.A(G2037_1003_gat), .Y(G2037_1003_ngat) );
INVXL U_g1933 (.A(G1984_1010_gat), .Y(G1984_1010_ngat) );
INVXL U_g1934 (.A(G1987_1004_gat), .Y(G1987_1004_ngat) );
INVXL U_g1935 (.A(G1883_1011_gat), .Y(G1883_1011_ngat) );
INVXL U_g1936 (.A(G1886_1005_gat), .Y(G1886_1005_ngat) );
INVXL U_g1937 (.A(G2254_993_gat), .Y(G2254_993_ngat) );
INVXL U_g1938 (.A(G2255_987_gat), .Y(G2255_987_ngat) );
INVXL U_g1939 (.A(G2256_959_gat), .Y(G2256_959_ngat) );
INVXL U_g1940 (.A(G2202_994_gat), .Y(G2202_994_ngat) );
INVXL U_g1941 (.A(G2203_988_gat), .Y(G2203_988_ngat) );
INVXL U_g1942 (.A(G2204_961_gat), .Y(G2204_961_ngat) );
INVXL U_g1943 (.A(G2111_1035_gat), .Y(G2111_1035_ngat) );
INVXL U_g1944 (.A(G2114_388_gat), .Y(G2114_388_ngat) );
INVXL U_g1945 (.A(G2117_531_gat), .Y(G2117_531_ngat) );
INVXL U_g1946 (.A(G2097_995_gat), .Y(G2097_995_ngat) );
INVXL U_g1947 (.A(G2098_989_gat), .Y(G2098_989_ngat) );
INVXL U_g1948 (.A(G2099_963_gat), .Y(G2099_963_ngat) );
INVXL U_g1949 (.A(G2040_996_gat), .Y(G2040_996_ngat) );
INVXL U_g1950 (.A(G2041_990_gat), .Y(G2041_990_ngat) );
INVXL U_g1951 (.A(G2042_964_gat), .Y(G2042_964_ngat) );
INVXL U_g1952 (.A(G1990_997_gat), .Y(G1990_997_ngat) );
INVXL U_g1953 (.A(G1991_991_gat), .Y(G1991_991_ngat) );
INVXL U_g1954 (.A(G1992_966_gat), .Y(G1992_966_ngat) );
INVXL U_g1955 (.A(G1903_1034_gat), .Y(G1903_1034_ngat) );
INVXL U_g1956 (.A(G1906_411_gat), .Y(G1906_411_ngat) );
INVXL U_g1957 (.A(G1909_545_gat), .Y(G1909_545_ngat) );
INVXL U_g1958 (.A(G1889_998_gat), .Y(G1889_998_ngat) );
INVXL U_g1959 (.A(G1890_992_gat), .Y(G1890_992_ngat) );
INVXL U_g1960 (.A(G1891_967_gat), .Y(G1891_967_ngat) );
INVXL U_g1961 (.A(G1536_1016_gat), .Y(G1536_1016_ngat) );
INVXL U_g1962 (.A(G1537_1018_gat), .Y(G1537_1018_ngat) );
INVXL U_g1963 (.A(G1538_548_gat), .Y(G1538_548_ngat) );
INVXL U_g1964 (.A(G679_1015_gat), .Y(G679_1015_ngat) );
INVXL U_g1965 (.A(G680_420_gat), .Y(G680_420_ngat) );
INVXL U_g1966 (.A(G669_1019_gat), .Y(G669_1019_ngat) );
INVXL U_g1967 (.A(G671_426_gat), .Y(G671_426_ngat) );
INVXL U_g1968 (.A(G672_533_gat), .Y(G672_533_ngat) );
INVXL U_g1969 (.A(G1582_1020_gat), .Y(G1582_1020_ngat) );
INVXL U_g1970 (.A(G1583_1021_gat), .Y(G1583_1021_ngat) );
INVXL U_g1971 (.A(G1586_1022_gat), .Y(G1586_1022_ngat) );
INVXL U_g1972 (.A(G1587_1023_gat), .Y(G1587_1023_ngat) );
INVXL U_g1973 (.A(G1590_1024_gat), .Y(G1590_1024_ngat) );
INVXL U_g1974 (.A(G1591_1025_gat), .Y(G1591_1025_ngat) );
INVXL U_g1975 (.A(G1594_1026_gat), .Y(G1594_1026_ngat) );
INVXL U_g1976 (.A(G1595_1027_gat), .Y(G1595_1027_ngat) );
INVXL U_g1977 (.A(G1598_1028_gat), .Y(G1598_1028_ngat) );
INVXL U_g1978 (.A(G1599_1029_gat), .Y(G1599_1029_ngat) );
INVXL U_g1979 (.A(G1602_1030_gat), .Y(G1602_1030_ngat) );
INVXL U_g1980 (.A(G1603_1031_gat), .Y(G1603_1031_ngat) );
INVXL U_g1981 (.A(G1606_1032_gat), .Y(G1606_1032_ngat) );
INVXL U_g1982 (.A(G1607_1033_gat), .Y(G1607_1033_ngat) );
INVXL U_g1983 (.A(G661_1080_gat), .Y(G661_1080_ngat) );
INVXL U_g1984 (.A(G662_550_gat), .Y(G662_550_ngat) );
INVXL U_g1985 (.A(G2149_1104_gat), .Y(G2149_1104_ngat) );
INVXL U_g1986 (.A(G2150_1102_gat), .Y(G2150_1102_ngat) );
INVXL U_g1987 (.A(G2151_1122_gat), .Y(G2151_1122_ngat) );
INVXL U_g1988 (.A(G1939_1105_gat), .Y(G1939_1105_ngat) );
INVXL U_g1989 (.A(G1940_1103_gat), .Y(G1940_1103_ngat) );
INVXL U_g1990 (.A(G1941_1123_gat), .Y(G1941_1123_ngat) );
INVXL U_g1991 (.A(G2143_1116_gat), .Y(G2143_1116_ngat) );
INVXL U_g1992 (.A(G2146_1108_gat), .Y(G2146_1108_ngat) );
INVXL U_g1993 (.A(G1933_1117_gat), .Y(G1933_1117_ngat) );
INVXL U_g1994 (.A(G1936_1113_gat), .Y(G1936_1113_ngat) );
INVXL U_g1995 (.A(G689_1125_gat), .Y(G689_1125_ngat) );
INVXL U_g1996 (.A(G690_535_gat), .Y(G690_535_ngat) );
INVXL U_g1997 (.A(G691_524_gat), .Y(G691_524_ngat) );
INVXL U_g1998 (.A(G700_1160_gat), .Y(G700_1160_ngat) );
INVXL U_g1999 (.A(G701_523_gat), .Y(G701_523_ngat) );
INVXL U_g2000 (.A(G702_530_gat), .Y(G702_530_ngat) );
INVXL U_g2001 (.A(G2489_1100_gat), .Y(G2489_1100_ngat) );
INVXL U_g2002 (.A(G2490_1230_gat), .Y(G2490_1230_ngat) );
INVXL U_g2003 (.A(G2455_1095_gat), .Y(G2455_1095_ngat) );
INVXL U_g2004 (.A(G2518_1274_gat), .Y(G2518_1274_ngat) );
INVXL U_g2005 (.A(G2448_1099_gat), .Y(G2448_1099_ngat) );
INVXL U_g2006 (.A(G2517_1302_gat), .Y(G2517_1302_ngat) );
INVXL U_g2007 (.A(G2275_1246_gat), .Y(G2275_1246_ngat) );
INVXL U_g2008 (.A(G2500_1319_gat), .Y(G2500_1319_ngat) );
INVXL U_g2009 (.A(G1639_1130_gat), .Y(G1639_1130_ngat) );
INVXL U_g2010 (.A(G1641_1327_gat), .Y(G1641_1327_ngat) );
INVXL U_g2011 (.A(G1643_727_gat), .Y(G1643_727_ngat) );
INVXL U_g2012 (.A(G1630_1129_gat), .Y(G1630_1129_ngat) );
INVXL U_g2013 (.A(G1632_1326_gat), .Y(G1632_1326_ngat) );
INVXL U_g2014 (.A(G1634_730_gat), .Y(G1634_730_ngat) );
INVXL U_g2015 (.A(G1612_1127_gat), .Y(G1612_1127_ngat) );
INVXL U_g2016 (.A(G1614_1325_gat), .Y(G1614_1325_ngat) );
INVXL U_g2017 (.A(G1616_733_gat), .Y(G1616_733_ngat) );
INVXL U_g2018 (.A(G1648_1131_gat), .Y(G1648_1131_ngat) );
INVXL U_g2019 (.A(G1650_1322_gat), .Y(G1650_1322_ngat) );
INVXL U_g2020 (.A(G1652_1090_gat), .Y(G1652_1090_ngat) );
INVXL U_g2021 (.A(G1666_1133_gat), .Y(G1666_1133_ngat) );
INVXL U_g2022 (.A(G1668_1323_gat), .Y(G1668_1323_ngat) );
INVXL U_g2023 (.A(G1670_1225_gat), .Y(G1670_1225_ngat) );
INVXL U_g2024 (.A(G1675_1134_gat), .Y(G1675_1134_ngat) );
INVXL U_g2025 (.A(G1677_1324_gat), .Y(G1677_1324_ngat) );
INVXL U_g2026 (.A(G1679_1188_gat), .Y(G1679_1188_ngat) );
INVXL U_g2027 (.A(G2643_1328_gat), .Y(G2643_1328_ngat) );
INVXL U_g2028 (.A(G2645_1305_gat), .Y(G2645_1305_ngat) );
INVXL U_g2029 (.A(G1621_1128_gat), .Y(G1621_1128_ngat) );
INVXL U_g2030 (.A(G1623_1387_gat), .Y(G1623_1387_ngat) );
INVXL U_g2031 (.A(G1625_732_gat), .Y(G1625_732_ngat) );
INVXL U_g2032 (.A(G1657_1132_gat), .Y(G1657_1132_ngat) );
INVXL U_g2033 (.A(G1659_1386_gat), .Y(G1659_1386_ngat) );
INVXL U_g2034 (.A(G1661_1126_gat), .Y(G1661_1126_ngat) );
INVXL U_g2035 (.A(G397_1394_gat), .Y(G397_1394_ngat) );
INVXL U_g2036 (.A(G398_1366_gat), .Y(G398_1366_ngat) );
INVXL U_g2037 (.A(G929_734_gat), .Y(G929_734_ngat) );
INVXL U_g2038 (.A(G933_1419_gat), .Y(G933_1419_ngat) );
INVXL U_g2039 (.A(G938_722_gat), .Y(G938_722_ngat) );
INVXL U_g2040 (.A(G2633_1420_gat), .Y(G2633_1420_ngat) );
INVXL U_g2041 (.A(G2634_1416_gat), .Y(G2634_1416_ngat) );
INVXL U_g2042 (.A(G2805_1446_gat), .Y(G2805_1446_ngat) );
INVXL U_g2043 (.A(G2808_1443_gat), .Y(G2808_1443_ngat) );
INVXL U_g2044 (.A(G2811_1393_gat), .Y(G2811_1393_ngat) );
INVXL U_g2045 (.A(G2736_1502_gat), .Y(G2736_1502_ngat) );
INVXL U_g2046 (.A(G2739_1501_gat), .Y(G2739_1501_ngat) );
INVXL U_g2047 (.A(G2742_1390_gat), .Y(G2742_1390_ngat) );
INVXL U_g2048 (.A(G2600_1542_gat), .Y(G2600_1542_ngat) );
INVXL U_g2049 (.A(G2650_1404_gat), .Y(G2650_1404_ngat) );
INVXL U_g2050 (.A(G2661_1561_gat), .Y(G2661_1561_ngat) );
INVXL U_g2051 (.A(G2662_1548_gat), .Y(G2662_1548_ngat) );
INVXL U_g2052 (.A(G944_969_gat), .Y(G944_969_ngat) );
INVXL U_g2053 (.A(G947_910_gat), .Y(G947_910_ngat) );
INVXL U_g2054 (.A(G951_1564_gat), .Y(G951_1564_ngat) );
INVXL U_g2055 (.A(G2555_1566_gat), .Y(G2555_1566_ngat) );
INVXL U_g2056 (.A(G2638_1483_gat), .Y(G2638_1483_ngat) );
INVXL U_g2057 (.A(G2771_1523_gat), .Y(G2771_1523_ngat) );
INVXL U_g2058 (.A(G2774_1572_gat), .Y(G2774_1572_ngat) );
INVXL U_g2059 (.A(G2777_1445_gat), .Y(G2777_1445_ngat) );
INVXL U_g2060 (.A(G2788_1503_gat), .Y(G2788_1503_ngat) );
INVXL U_g2061 (.A(G2791_1573_gat), .Y(G2791_1573_ngat) );
INVXL U_g2062 (.A(G2794_1392_gat), .Y(G2794_1392_ngat) );
INVXL U_g2063 (.A(G2658_1575_gat), .Y(G2658_1575_ngat) );
INVXL U_g2064 (.A(G2659_1568_gat), .Y(G2659_1568_ngat) );
INVXL U_g2065 (.A(G2700_1520_gat), .Y(G2700_1520_ngat) );
INVXL U_g2066 (.A(G2703_1578_gat), .Y(G2703_1578_ngat) );
INVXL U_g2067 (.A(G2706_1444_gat), .Y(G2706_1444_ngat) );
INVXL U_g2068 (.A(G2754_1556_gat), .Y(G2754_1556_ngat) );
INVXL U_g2069 (.A(G2757_1579_gat), .Y(G2757_1579_ngat) );
INVXL U_g2070 (.A(G2760_1391_gat), .Y(G2760_1391_ngat) );
INVXL U_g2071 (.A(G2719_1538_gat), .Y(G2719_1538_ngat) );
INVXL U_g2072 (.A(G2722_1586_gat), .Y(G2722_1586_ngat) );
INVXL U_g2073 (.A(G2725_1389_gat), .Y(G2725_1389_ngat) );
INVXL U_g2074 (.A(G2681_1574_gat), .Y(G2681_1574_ngat) );
INVXL U_g2075 (.A(G2684_1596_gat), .Y(G2684_1596_ngat) );
INVXL U_g2076 (.A(G2687_1388_gat), .Y(G2687_1388_ngat) );
INVXL U_g2077 (.A(G2928_1623_gat), .Y(G2928_1623_ngat) );
INVXL U_g2078 (.A(G2929_1644_gat), .Y(G2929_1644_ngat) );
INVXL U_g2079 (.A(G2906_1677_gat), .Y(G2906_1677_ngat) );
INVXL U_g2080 (.A(G2907_1683_gat), .Y(G2907_1683_ngat) );
INVXL U_g2081 (.A(G2908_1676_gat), .Y(G2908_1676_ngat) );
INVXL U_g2082 (.A(G2909_1684_gat), .Y(G2909_1684_ngat) );

endmodule
