module C499 ( GID0_0_gat, GID1_1_gat, GID2_2_gat, GID3_3_gat, GID4_4_gat, GID5_5_gat, GID6_6_gat, GID7_7_gat, GID8_8_gat, GID9_9_gat, GID10_10_gat, GID11_11_gat, GID12_12_gat, GID13_13_gat, GID14_14_gat, GID15_15_gat, GID16_16_gat, GID17_17_gat, GID18_18_gat, GID19_19_gat, GID20_20_gat, GID21_21_gat, GID22_22_gat, GID23_23_gat, GID24_24_gat, GID25_25_gat, GID26_26_gat, GID27_27_gat, GID28_28_gat, GID29_29_gat, GID30_30_gat, GID31_31_gat, GIC0_32_gat, GIC1_33_gat, GIC2_34_gat, GIC3_35_gat, GIC4_36_gat, GIC5_37_gat, GIC6_38_gat, GIC7_39_gat, GR_40_gat, GOD0_242_gat, GOD1_241_gat, GOD2_240_gat, GOD3_239_gat, GOD4_238_gat, GOD5_237_gat, GOD6_236_gat, GOD7_235_gat, GOD8_234_gat, GOD9_233_gat, GOD10_232_gat, GOD11_231_gat, GOD12_230_gat, GOD13_229_gat, GOD14_228_gat, GOD15_227_gat, GOD16_226_gat, GOD17_225_gat, GOD18_224_gat, GOD19_223_gat, GOD20_222_gat, GOD21_221_gat, GOD22_220_gat, GOD23_219_gat, GOD24_218_gat, GOD25_217_gat, GOD26_216_gat, GOD27_215_gat, GOD28_214_gat, GOD29_213_gat, GOD30_212_gat, GOD31_211_gat);

input GID0_0_gat;
input GID1_1_gat;
input GID2_2_gat;
input GID3_3_gat;
input GID4_4_gat;
input GID5_5_gat;
input GID6_6_gat;
input GID7_7_gat;
input GID8_8_gat;
input GID9_9_gat;
input GID10_10_gat;
input GID11_11_gat;
input GID12_12_gat;
input GID13_13_gat;
input GID14_14_gat;
input GID15_15_gat;
input GID16_16_gat;
input GID17_17_gat;
input GID18_18_gat;
input GID19_19_gat;
input GID20_20_gat;
input GID21_21_gat;
input GID22_22_gat;
input GID23_23_gat;
input GID24_24_gat;
input GID25_25_gat;
input GID26_26_gat;
input GID27_27_gat;
input GID28_28_gat;
input GID29_29_gat;
input GID30_30_gat;
input GID31_31_gat;
input GIC0_32_gat;
input GIC1_33_gat;
input GIC2_34_gat;
input GIC3_35_gat;
input GIC4_36_gat;
input GIC5_37_gat;
input GIC6_38_gat;
input GIC7_39_gat;
input GR_40_gat;

output GOD0_242_gat;
output GOD1_241_gat;
output GOD2_240_gat;
output GOD3_239_gat;
output GOD4_238_gat;
output GOD5_237_gat;
output GOD6_236_gat;
output GOD7_235_gat;
output GOD8_234_gat;
output GOD9_233_gat;
output GOD10_232_gat;
output GOD11_231_gat;
output GOD12_230_gat;
output GOD13_229_gat;
output GOD14_228_gat;
output GOD15_227_gat;
output GOD16_226_gat;
output GOD17_225_gat;
output GOD18_224_gat;
output GOD19_223_gat;
output GOD20_222_gat;
output GOD21_221_gat;
output GOD22_220_gat;
output GOD23_219_gat;
output GOD24_218_gat;
output GOD25_217_gat;
output GOD26_216_gat;
output GOD27_215_gat;
output GOD28_214_gat;
output GOD29_213_gat;
output GOD30_212_gat;
output GOD31_211_gat;

AND2XL U_g1 (.A(GR_40_gat), .B(GIC7_39_gat), .Y(GH7_41_gat) );
AND2XL U_g2 (.A(GR_40_gat), .B(GIC6_38_gat), .Y(GH6_42_gat) );
AND2XL U_g3 (.A(GR_40_gat), .B(GIC5_37_gat), .Y(GH5_43_gat) );
AND2XL U_g4 (.A(GR_40_gat), .B(GIC4_36_gat), .Y(GH4_44_gat) );
AND2XL U_g5 (.A(GR_40_gat), .B(GIC3_35_gat), .Y(GH3_45_gat) );
AND2XL U_g6 (.A(GR_40_gat), .B(GIC2_34_gat), .Y(GH2_46_gat) );
AND2XL U_g7 (.A(GR_40_gat), .B(GIC1_33_gat), .Y(GH1_47_gat) );
AND2XL U_g8 (.A(GR_40_gat), .B(GIC0_32_gat), .Y(GH0_48_gat) );
OR2XL U_g9 (.A(Ginternal__11gat), .B(Ginternal__10gat), .Y(GXA15_49_gat) );
AND2XL U_g10 (.A(GID31_31_gat), .B(GID30_30_ngat), .Y(Ginternal__10gat) );
AND2XL U_g11 (.A(GID31_31_ngat), .B(GID30_30_gat), .Y(Ginternal__11gat) );
OR2XL U_g12 (.A(Ginternal__14gat), .B(Ginternal__13gat), .Y(GXA14_50_gat) );
AND2XL U_g13 (.A(GID29_29_gat), .B(GID28_28_ngat), .Y(Ginternal__13gat) );
AND2XL U_g14 (.A(GID29_29_ngat), .B(GID28_28_gat), .Y(Ginternal__14gat) );
OR2XL U_g15 (.A(Ginternal__17gat), .B(Ginternal__16gat), .Y(GXC7_51_gat) );
AND2XL U_g16 (.A(GID31_31_gat), .B(GID27_27_ngat), .Y(Ginternal__16gat) );
AND2XL U_g17 (.A(GID31_31_ngat), .B(GID27_27_gat), .Y(Ginternal__17gat) );
OR2XL U_g18 (.A(Ginternal__20gat), .B(Ginternal__19gat), .Y(GXC6_52_gat) );
AND2XL U_g19 (.A(GID30_30_gat), .B(GID26_26_ngat), .Y(Ginternal__19gat) );
AND2XL U_g20 (.A(GID30_30_ngat), .B(GID26_26_gat), .Y(Ginternal__20gat) );
OR2XL U_g21 (.A(Ginternal__23gat), .B(Ginternal__22gat), .Y(GXA13_53_gat) );
AND2XL U_g22 (.A(GID27_27_gat), .B(GID26_26_ngat), .Y(Ginternal__22gat) );
AND2XL U_g23 (.A(GID27_27_ngat), .B(GID26_26_gat), .Y(Ginternal__23gat) );
OR2XL U_g24 (.A(Ginternal__26gat), .B(Ginternal__25gat), .Y(GXC5_54_gat) );
AND2XL U_g25 (.A(GID29_29_gat), .B(GID25_25_ngat), .Y(Ginternal__25gat) );
AND2XL U_g26 (.A(GID29_29_ngat), .B(GID25_25_gat), .Y(Ginternal__26gat) );
OR2XL U_g27 (.A(Ginternal__29gat), .B(Ginternal__28gat), .Y(GXC4_55_gat) );
AND2XL U_g28 (.A(GID28_28_gat), .B(GID24_24_ngat), .Y(Ginternal__28gat) );
AND2XL U_g29 (.A(GID28_28_ngat), .B(GID24_24_gat), .Y(Ginternal__29gat) );
OR2XL U_g30 (.A(Ginternal__32gat), .B(Ginternal__31gat), .Y(GXA12_56_gat) );
AND2XL U_g31 (.A(GID25_25_gat), .B(GID24_24_ngat), .Y(Ginternal__31gat) );
AND2XL U_g32 (.A(GID25_25_ngat), .B(GID24_24_gat), .Y(Ginternal__32gat) );
OR2XL U_g33 (.A(Ginternal__35gat), .B(Ginternal__34gat), .Y(GXA11_57_gat) );
AND2XL U_g34 (.A(GID23_23_gat), .B(GID22_22_ngat), .Y(Ginternal__34gat) );
AND2XL U_g35 (.A(GID23_23_ngat), .B(GID22_22_gat), .Y(Ginternal__35gat) );
OR2XL U_g36 (.A(Ginternal__38gat), .B(Ginternal__37gat), .Y(GXA10_58_gat) );
AND2XL U_g37 (.A(GID21_21_gat), .B(GID20_20_ngat), .Y(Ginternal__37gat) );
AND2XL U_g38 (.A(GID21_21_ngat), .B(GID20_20_gat), .Y(Ginternal__38gat) );
OR2XL U_g39 (.A(Ginternal__41gat), .B(Ginternal__40gat), .Y(GXB7_59_gat) );
AND2XL U_g40 (.A(GID23_23_gat), .B(GID19_19_ngat), .Y(Ginternal__40gat) );
AND2XL U_g41 (.A(GID23_23_ngat), .B(GID19_19_gat), .Y(Ginternal__41gat) );
OR2XL U_g42 (.A(Ginternal__44gat), .B(Ginternal__43gat), .Y(GXB6_60_gat) );
AND2XL U_g43 (.A(GID22_22_gat), .B(GID18_18_ngat), .Y(Ginternal__43gat) );
AND2XL U_g44 (.A(GID22_22_ngat), .B(GID18_18_gat), .Y(Ginternal__44gat) );
OR2XL U_g45 (.A(Ginternal__47gat), .B(Ginternal__46gat), .Y(GXA9_61_gat) );
AND2XL U_g46 (.A(GID19_19_gat), .B(GID18_18_ngat), .Y(Ginternal__46gat) );
AND2XL U_g47 (.A(GID19_19_ngat), .B(GID18_18_gat), .Y(Ginternal__47gat) );
OR2XL U_g48 (.A(Ginternal__50gat), .B(Ginternal__49gat), .Y(GXB5_62_gat) );
AND2XL U_g49 (.A(GID21_21_gat), .B(GID17_17_ngat), .Y(Ginternal__49gat) );
AND2XL U_g50 (.A(GID21_21_ngat), .B(GID17_17_gat), .Y(Ginternal__50gat) );
OR2XL U_g51 (.A(Ginternal__53gat), .B(Ginternal__52gat), .Y(GXB4_63_gat) );
AND2XL U_g52 (.A(GID20_20_gat), .B(GID16_16_ngat), .Y(Ginternal__52gat) );
AND2XL U_g53 (.A(GID20_20_ngat), .B(GID16_16_gat), .Y(Ginternal__53gat) );
OR2XL U_g54 (.A(Ginternal__56gat), .B(Ginternal__55gat), .Y(GXA8_64_gat) );
AND2XL U_g55 (.A(GID17_17_gat), .B(GID16_16_ngat), .Y(Ginternal__55gat) );
AND2XL U_g56 (.A(GID17_17_ngat), .B(GID16_16_gat), .Y(Ginternal__56gat) );
OR2XL U_g57 (.A(Ginternal__59gat), .B(Ginternal__58gat), .Y(GXA7_65_gat) );
AND2XL U_g58 (.A(GID15_15_gat), .B(GID14_14_ngat), .Y(Ginternal__58gat) );
AND2XL U_g59 (.A(GID15_15_ngat), .B(GID14_14_gat), .Y(Ginternal__59gat) );
OR2XL U_g60 (.A(Ginternal__62gat), .B(Ginternal__61gat), .Y(GXA6_66_gat) );
AND2XL U_g61 (.A(GID13_13_gat), .B(GID12_12_ngat), .Y(Ginternal__61gat) );
AND2XL U_g62 (.A(GID13_13_ngat), .B(GID12_12_gat), .Y(Ginternal__62gat) );
OR2XL U_g63 (.A(Ginternal__65gat), .B(Ginternal__64gat), .Y(GXC3_67_gat) );
AND2XL U_g64 (.A(GID15_15_gat), .B(GID11_11_ngat), .Y(Ginternal__64gat) );
AND2XL U_g65 (.A(GID15_15_ngat), .B(GID11_11_gat), .Y(Ginternal__65gat) );
OR2XL U_g66 (.A(Ginternal__68gat), .B(Ginternal__67gat), .Y(GXC2_68_gat) );
AND2XL U_g67 (.A(GID14_14_gat), .B(GID10_10_ngat), .Y(Ginternal__67gat) );
AND2XL U_g68 (.A(GID14_14_ngat), .B(GID10_10_gat), .Y(Ginternal__68gat) );
OR2XL U_g69 (.A(Ginternal__71gat), .B(Ginternal__70gat), .Y(GXA5_69_gat) );
AND2XL U_g70 (.A(GID11_11_gat), .B(GID10_10_ngat), .Y(Ginternal__70gat) );
AND2XL U_g71 (.A(GID11_11_ngat), .B(GID10_10_gat), .Y(Ginternal__71gat) );
OR2XL U_g72 (.A(Ginternal__74gat), .B(Ginternal__73gat), .Y(GXC1_70_gat) );
AND2XL U_g73 (.A(GID13_13_gat), .B(GID9_9_ngat), .Y(Ginternal__73gat) );
AND2XL U_g74 (.A(GID13_13_ngat), .B(GID9_9_gat), .Y(Ginternal__74gat) );
OR2XL U_g75 (.A(Ginternal__77gat), .B(Ginternal__76gat), .Y(GXC0_71_gat) );
AND2XL U_g76 (.A(GID12_12_gat), .B(GID8_8_ngat), .Y(Ginternal__76gat) );
AND2XL U_g77 (.A(GID12_12_ngat), .B(GID8_8_gat), .Y(Ginternal__77gat) );
OR2XL U_g78 (.A(Ginternal__80gat), .B(Ginternal__79gat), .Y(GXA4_72_gat) );
AND2XL U_g79 (.A(GID9_9_gat), .B(GID8_8_ngat), .Y(Ginternal__79gat) );
AND2XL U_g80 (.A(GID9_9_ngat), .B(GID8_8_gat), .Y(Ginternal__80gat) );
OR2XL U_g81 (.A(Ginternal__83gat), .B(Ginternal__82gat), .Y(GXA3_73_gat) );
AND2XL U_g82 (.A(GID7_7_gat), .B(GID6_6_ngat), .Y(Ginternal__82gat) );
AND2XL U_g83 (.A(GID7_7_ngat), .B(GID6_6_gat), .Y(Ginternal__83gat) );
OR2XL U_g84 (.A(Ginternal__86gat), .B(Ginternal__85gat), .Y(GXA2_74_gat) );
AND2XL U_g85 (.A(GID5_5_gat), .B(GID4_4_ngat), .Y(Ginternal__85gat) );
AND2XL U_g86 (.A(GID5_5_ngat), .B(GID4_4_gat), .Y(Ginternal__86gat) );
OR2XL U_g87 (.A(Ginternal__89gat), .B(Ginternal__88gat), .Y(GXB3_75_gat) );
AND2XL U_g88 (.A(GID7_7_gat), .B(GID3_3_ngat), .Y(Ginternal__88gat) );
AND2XL U_g89 (.A(GID7_7_ngat), .B(GID3_3_gat), .Y(Ginternal__89gat) );
OR2XL U_g90 (.A(Ginternal__92gat), .B(Ginternal__91gat), .Y(GXB2_76_gat) );
AND2XL U_g91 (.A(GID6_6_gat), .B(GID2_2_ngat), .Y(Ginternal__91gat) );
AND2XL U_g92 (.A(GID6_6_ngat), .B(GID2_2_gat), .Y(Ginternal__92gat) );
OR2XL U_g93 (.A(Ginternal__95gat), .B(Ginternal__94gat), .Y(GXA1_77_gat) );
AND2XL U_g94 (.A(GID3_3_gat), .B(GID2_2_ngat), .Y(Ginternal__94gat) );
AND2XL U_g95 (.A(GID3_3_ngat), .B(GID2_2_gat), .Y(Ginternal__95gat) );
OR2XL U_g96 (.A(Ginternal__98gat), .B(Ginternal__97gat), .Y(GXB1_78_gat) );
AND2XL U_g97 (.A(GID5_5_gat), .B(GID1_1_ngat), .Y(Ginternal__97gat) );
AND2XL U_g98 (.A(GID5_5_ngat), .B(GID1_1_gat), .Y(Ginternal__98gat) );
OR2XL U_g99 (.A(Ginternal__101gat), .B(Ginternal__100gat), .Y(GXB0_79_gat) );
AND2XL U_g100 (.A(GID4_4_gat), .B(GID0_0_ngat), .Y(Ginternal__100gat) );
AND2XL U_g101 (.A(GID4_4_ngat), .B(GID0_0_gat), .Y(Ginternal__101gat) );
OR2XL U_g102 (.A(Ginternal__104gat), .B(Ginternal__103gat), .Y(GXA0_80_gat) );
AND2XL U_g103 (.A(GID1_1_gat), .B(GID0_0_ngat), .Y(Ginternal__103gat) );
AND2XL U_g104 (.A(GID1_1_ngat), .B(GID0_0_gat), .Y(Ginternal__104gat) );
OR2XL U_g105 (.A(Ginternal__107gat), .B(Ginternal__106gat), .Y(GF7_81_gat) );
AND2XL U_g106 (.A(GXA15_49_gat), .B(GXA14_50_ngat), .Y(Ginternal__106gat) );
AND2XL U_g107 (.A(GXA15_49_ngat), .B(GXA14_50_gat), .Y(Ginternal__107gat) );
OR2XL U_g108 (.A(Ginternal__110gat), .B(Ginternal__109gat), .Y(GXE7_82_gat) );
AND2XL U_g109 (.A(GXC7_51_gat), .B(GXB7_59_ngat), .Y(Ginternal__109gat) );
AND2XL U_g110 (.A(GXC7_51_ngat), .B(GXB7_59_gat), .Y(Ginternal__110gat) );
OR2XL U_g111 (.A(Ginternal__113gat), .B(Ginternal__112gat), .Y(GXE6_83_gat) );
AND2XL U_g112 (.A(GXC6_52_gat), .B(GXB6_60_ngat), .Y(Ginternal__112gat) );
AND2XL U_g113 (.A(GXC6_52_ngat), .B(GXB6_60_gat), .Y(Ginternal__113gat) );
OR2XL U_g114 (.A(Ginternal__116gat), .B(Ginternal__115gat), .Y(GF6_84_gat) );
AND2XL U_g115 (.A(GXA13_53_gat), .B(GXA12_56_ngat), .Y(Ginternal__115gat) );
AND2XL U_g116 (.A(GXA13_53_ngat), .B(GXA12_56_gat), .Y(Ginternal__116gat) );
OR2XL U_g117 (.A(Ginternal__119gat), .B(Ginternal__118gat), .Y(GXE5_85_gat) );
AND2XL U_g118 (.A(GXC5_54_gat), .B(GXB5_62_ngat), .Y(Ginternal__118gat) );
AND2XL U_g119 (.A(GXC5_54_ngat), .B(GXB5_62_gat), .Y(Ginternal__119gat) );
OR2XL U_g120 (.A(Ginternal__122gat), .B(Ginternal__121gat), .Y(GXE4_86_gat) );
AND2XL U_g121 (.A(GXC4_55_gat), .B(GXB4_63_ngat), .Y(Ginternal__121gat) );
AND2XL U_g122 (.A(GXC4_55_ngat), .B(GXB4_63_gat), .Y(Ginternal__122gat) );
OR2XL U_g123 (.A(Ginternal__125gat), .B(Ginternal__124gat), .Y(GF5_87_gat) );
AND2XL U_g124 (.A(GXA11_57_gat), .B(GXA10_58_ngat), .Y(Ginternal__124gat) );
AND2XL U_g125 (.A(GXA11_57_ngat), .B(GXA10_58_gat), .Y(Ginternal__125gat) );
OR2XL U_g126 (.A(Ginternal__128gat), .B(Ginternal__127gat), .Y(GF4_88_gat) );
AND2XL U_g127 (.A(GXA9_61_gat), .B(GXA8_64_ngat), .Y(Ginternal__127gat) );
AND2XL U_g128 (.A(GXA9_61_ngat), .B(GXA8_64_gat), .Y(Ginternal__128gat) );
OR2XL U_g129 (.A(Ginternal__131gat), .B(Ginternal__130gat), .Y(GF3_89_gat) );
AND2XL U_g130 (.A(GXA7_65_gat), .B(GXA6_66_ngat), .Y(Ginternal__130gat) );
AND2XL U_g131 (.A(GXA7_65_ngat), .B(GXA6_66_gat), .Y(Ginternal__131gat) );
OR2XL U_g132 (.A(Ginternal__134gat), .B(Ginternal__133gat), .Y(GXE3_90_gat) );
AND2XL U_g133 (.A(GXC3_67_gat), .B(GXB3_75_ngat), .Y(Ginternal__133gat) );
AND2XL U_g134 (.A(GXC3_67_ngat), .B(GXB3_75_gat), .Y(Ginternal__134gat) );
OR2XL U_g135 (.A(Ginternal__137gat), .B(Ginternal__136gat), .Y(GXE2_91_gat) );
AND2XL U_g136 (.A(GXC2_68_gat), .B(GXB2_76_ngat), .Y(Ginternal__136gat) );
AND2XL U_g137 (.A(GXC2_68_ngat), .B(GXB2_76_gat), .Y(Ginternal__137gat) );
OR2XL U_g138 (.A(Ginternal__140gat), .B(Ginternal__139gat), .Y(GF2_92_gat) );
AND2XL U_g139 (.A(GXA5_69_gat), .B(GXA4_72_ngat), .Y(Ginternal__139gat) );
AND2XL U_g140 (.A(GXA5_69_ngat), .B(GXA4_72_gat), .Y(Ginternal__140gat) );
OR2XL U_g141 (.A(Ginternal__143gat), .B(Ginternal__142gat), .Y(GXE1_93_gat) );
AND2XL U_g142 (.A(GXC1_70_gat), .B(GXB1_78_ngat), .Y(Ginternal__142gat) );
AND2XL U_g143 (.A(GXC1_70_ngat), .B(GXB1_78_gat), .Y(Ginternal__143gat) );
OR2XL U_g144 (.A(Ginternal__146gat), .B(Ginternal__145gat), .Y(GXE0_94_gat) );
AND2XL U_g145 (.A(GXC0_71_gat), .B(GXB0_79_ngat), .Y(Ginternal__145gat) );
AND2XL U_g146 (.A(GXC0_71_ngat), .B(GXB0_79_gat), .Y(Ginternal__146gat) );
OR2XL U_g147 (.A(Ginternal__149gat), .B(Ginternal__148gat), .Y(GF1_95_gat) );
AND2XL U_g148 (.A(GXA3_73_gat), .B(GXA2_74_ngat), .Y(Ginternal__148gat) );
AND2XL U_g149 (.A(GXA3_73_ngat), .B(GXA2_74_gat), .Y(Ginternal__149gat) );
OR2XL U_g150 (.A(Ginternal__152gat), .B(Ginternal__151gat), .Y(GF0_96_gat) );
AND2XL U_g151 (.A(GXA1_77_gat), .B(GXA0_80_ngat), .Y(Ginternal__151gat) );
AND2XL U_g152 (.A(GXA1_77_ngat), .B(GXA0_80_gat), .Y(Ginternal__152gat) );
OR2XL U_g153 (.A(Ginternal__155gat), .B(Ginternal__154gat), .Y(GG5_97_gat) );
AND2XL U_g154 (.A(GF7_81_gat), .B(GF6_84_ngat), .Y(Ginternal__154gat) );
AND2XL U_g155 (.A(GF7_81_ngat), .B(GF6_84_gat), .Y(Ginternal__155gat) );
OR2XL U_g156 (.A(Ginternal__158gat), .B(Ginternal__157gat), .Y(GG7_98_gat) );
AND2XL U_g157 (.A(GF7_81_gat), .B(GF5_87_ngat), .Y(Ginternal__157gat) );
AND2XL U_g158 (.A(GF7_81_ngat), .B(GF5_87_gat), .Y(Ginternal__158gat) );
OR2XL U_g159 (.A(Ginternal__161gat), .B(Ginternal__160gat), .Y(GG6_99_gat) );
AND2XL U_g160 (.A(GF6_84_gat), .B(GF4_88_ngat), .Y(Ginternal__160gat) );
AND2XL U_g161 (.A(GF6_84_ngat), .B(GF4_88_gat), .Y(Ginternal__161gat) );
OR2XL U_g162 (.A(Ginternal__164gat), .B(Ginternal__163gat), .Y(GG4_100_gat) );
AND2XL U_g163 (.A(GF5_87_gat), .B(GF4_88_ngat), .Y(Ginternal__163gat) );
AND2XL U_g164 (.A(GF5_87_ngat), .B(GF4_88_gat), .Y(Ginternal__164gat) );
OR2XL U_g165 (.A(Ginternal__167gat), .B(Ginternal__166gat), .Y(GG1_101_gat) );
AND2XL U_g166 (.A(GF3_89_gat), .B(GF2_92_ngat), .Y(Ginternal__166gat) );
AND2XL U_g167 (.A(GF3_89_ngat), .B(GF2_92_gat), .Y(Ginternal__167gat) );
OR2XL U_g168 (.A(Ginternal__170gat), .B(Ginternal__169gat), .Y(GG3_102_gat) );
AND2XL U_g169 (.A(GF3_89_gat), .B(GF1_95_ngat), .Y(Ginternal__169gat) );
AND2XL U_g170 (.A(GF3_89_ngat), .B(GF1_95_gat), .Y(Ginternal__170gat) );
OR2XL U_g171 (.A(Ginternal__173gat), .B(Ginternal__172gat), .Y(GG2_103_gat) );
AND2XL U_g172 (.A(GF2_92_gat), .B(GF0_96_ngat), .Y(Ginternal__172gat) );
AND2XL U_g173 (.A(GF2_92_ngat), .B(GF0_96_gat), .Y(Ginternal__173gat) );
OR2XL U_g174 (.A(Ginternal__176gat), .B(Ginternal__175gat), .Y(GG0_104_gat) );
AND2XL U_g175 (.A(GF1_95_gat), .B(GF0_96_ngat), .Y(Ginternal__175gat) );
AND2XL U_g176 (.A(GF1_95_ngat), .B(GF0_96_gat), .Y(Ginternal__176gat) );
OR2XL U_g177 (.A(Ginternal__179gat), .B(Ginternal__178gat), .Y(GXD7_105_gat) );
AND2XL U_g178 (.A(GG3_102_gat), .B(GH7_41_ngat), .Y(Ginternal__178gat) );
AND2XL U_g179 (.A(GG3_102_ngat), .B(GH7_41_gat), .Y(Ginternal__179gat) );
OR2XL U_g180 (.A(Ginternal__182gat), .B(Ginternal__181gat), .Y(GXD6_106_gat) );
AND2XL U_g181 (.A(GG2_103_gat), .B(GH6_42_ngat), .Y(Ginternal__181gat) );
AND2XL U_g182 (.A(GG2_103_ngat), .B(GH6_42_gat), .Y(Ginternal__182gat) );
OR2XL U_g183 (.A(Ginternal__185gat), .B(Ginternal__184gat), .Y(GXD5_107_gat) );
AND2XL U_g184 (.A(GG1_101_gat), .B(GH5_43_ngat), .Y(Ginternal__184gat) );
AND2XL U_g185 (.A(GG1_101_ngat), .B(GH5_43_gat), .Y(Ginternal__185gat) );
OR2XL U_g186 (.A(Ginternal__188gat), .B(Ginternal__187gat), .Y(GXD4_108_gat) );
AND2XL U_g187 (.A(GG0_104_gat), .B(GH4_44_ngat), .Y(Ginternal__187gat) );
AND2XL U_g188 (.A(GG0_104_ngat), .B(GH4_44_gat), .Y(Ginternal__188gat) );
OR2XL U_g189 (.A(Ginternal__191gat), .B(Ginternal__190gat), .Y(GXD3_109_gat) );
AND2XL U_g190 (.A(GG7_98_gat), .B(GH3_45_ngat), .Y(Ginternal__190gat) );
AND2XL U_g191 (.A(GG7_98_ngat), .B(GH3_45_gat), .Y(Ginternal__191gat) );
OR2XL U_g192 (.A(Ginternal__194gat), .B(Ginternal__193gat), .Y(GXD2_110_gat) );
AND2XL U_g193 (.A(GG6_99_gat), .B(GH2_46_ngat), .Y(Ginternal__193gat) );
AND2XL U_g194 (.A(GG6_99_ngat), .B(GH2_46_gat), .Y(Ginternal__194gat) );
OR2XL U_g195 (.A(Ginternal__197gat), .B(Ginternal__196gat), .Y(GXD1_111_gat) );
AND2XL U_g196 (.A(GG5_97_gat), .B(GH1_47_ngat), .Y(Ginternal__196gat) );
AND2XL U_g197 (.A(GG5_97_ngat), .B(GH1_47_gat), .Y(Ginternal__197gat) );
OR2XL U_g198 (.A(Ginternal__200gat), .B(Ginternal__199gat), .Y(GXD0_112_gat) );
AND2XL U_g199 (.A(GG4_100_gat), .B(GH0_48_ngat), .Y(Ginternal__199gat) );
AND2XL U_g200 (.A(GG4_100_ngat), .B(GH0_48_gat), .Y(Ginternal__200gat) );
OR2XL U_g201 (.A(Ginternal__203gat), .B(Ginternal__202gat), .Y(GS7_113_gat) );
AND2XL U_g202 (.A(GXD7_105_gat), .B(GXE7_82_ngat), .Y(Ginternal__202gat) );
AND2XL U_g203 (.A(GXD7_105_ngat), .B(GXE7_82_gat), .Y(Ginternal__203gat) );
OR2XL U_g204 (.A(Ginternal__206gat), .B(Ginternal__205gat), .Y(GS6_114_gat) );
AND2XL U_g205 (.A(GXD6_106_gat), .B(GXE6_83_ngat), .Y(Ginternal__205gat) );
AND2XL U_g206 (.A(GXD6_106_ngat), .B(GXE6_83_gat), .Y(Ginternal__206gat) );
OR2XL U_g207 (.A(Ginternal__209gat), .B(Ginternal__208gat), .Y(GS5_115_gat) );
AND2XL U_g208 (.A(GXD5_107_gat), .B(GXE5_85_ngat), .Y(Ginternal__208gat) );
AND2XL U_g209 (.A(GXD5_107_ngat), .B(GXE5_85_gat), .Y(Ginternal__209gat) );
OR2XL U_g210 (.A(Ginternal__212gat), .B(Ginternal__211gat), .Y(GS4_116_gat) );
AND2XL U_g211 (.A(GXD4_108_gat), .B(GXE4_86_ngat), .Y(Ginternal__211gat) );
AND2XL U_g212 (.A(GXD4_108_ngat), .B(GXE4_86_gat), .Y(Ginternal__212gat) );
OR2XL U_g213 (.A(Ginternal__215gat), .B(Ginternal__214gat), .Y(GS3_117_gat) );
AND2XL U_g214 (.A(GXD3_109_gat), .B(GXE3_90_ngat), .Y(Ginternal__214gat) );
AND2XL U_g215 (.A(GXD3_109_ngat), .B(GXE3_90_gat), .Y(Ginternal__215gat) );
OR2XL U_g216 (.A(Ginternal__218gat), .B(Ginternal__217gat), .Y(GS2_118_gat) );
AND2XL U_g217 (.A(GXD2_110_gat), .B(GXE2_91_ngat), .Y(Ginternal__217gat) );
AND2XL U_g218 (.A(GXD2_110_ngat), .B(GXE2_91_gat), .Y(Ginternal__218gat) );
OR2XL U_g219 (.A(Ginternal__221gat), .B(Ginternal__220gat), .Y(GS1_119_gat) );
AND2XL U_g220 (.A(GXD1_111_gat), .B(GXE1_93_ngat), .Y(Ginternal__220gat) );
AND2XL U_g221 (.A(GXD1_111_ngat), .B(GXE1_93_gat), .Y(Ginternal__221gat) );
OR2XL U_g222 (.A(Ginternal__224gat), .B(Ginternal__223gat), .Y(GS0_120_gat) );
AND2XL U_g223 (.A(GXD0_112_gat), .B(GXE0_94_ngat), .Y(Ginternal__223gat) );
AND2XL U_g224 (.A(GXD0_112_ngat), .B(GXE0_94_gat), .Y(Ginternal__224gat) );
BUFX20 U_g225 (.A(GS7_113_gat), .Y(GY7B_121_gat) );
BUFX20 U_g226 (.A(GS7_113_gat), .Y(GY7C_122_gat) );
BUFX20 U_g227 (.A(GS7_113_gat), .Y(GY7D_123_gat) );
BUFX20 U_g228 (.A(GS7_113_gat), .Y(GY7I_124_gat) );
BUFX20 U_g229 (.A(GS7_113_gat), .Y(GY7K_125_gat) );
BUFX20 U_g230 (.A(GS6_114_gat), .Y(GY6A_126_gat) );
BUFX20 U_g231 (.A(GS6_114_gat), .Y(GY6C_127_gat) );
BUFX20 U_g232 (.A(GS6_114_gat), .Y(GY6D_128_gat) );
BUFX20 U_g233 (.A(GS6_114_gat), .Y(GY6J_129_gat) );
BUFX20 U_g234 (.A(GS6_114_gat), .Y(GY6L_130_gat) );
BUFX20 U_g235 (.A(GS5_115_gat), .Y(GY5A_131_gat) );
BUFX20 U_g236 (.A(GS5_115_gat), .Y(GY5B_132_gat) );
BUFX20 U_g237 (.A(GS5_115_gat), .Y(GY5D_133_gat) );
BUFX20 U_g238 (.A(GS5_115_gat), .Y(GY5I_134_gat) );
BUFX20 U_g239 (.A(GS5_115_gat), .Y(GY5J_135_gat) );
BUFX20 U_g240 (.A(GS4_116_gat), .Y(GY4A_136_gat) );
BUFX20 U_g241 (.A(GS4_116_gat), .Y(GY4B_137_gat) );
BUFX20 U_g242 (.A(GS4_116_gat), .Y(GY4C_138_gat) );
BUFX20 U_g243 (.A(GS4_116_gat), .Y(GY4K_139_gat) );
BUFX20 U_g244 (.A(GS4_116_gat), .Y(GY4L_140_gat) );
BUFX20 U_g245 (.A(GS3_117_gat), .Y(GY3B_141_gat) );
BUFX20 U_g246 (.A(GS3_117_gat), .Y(GY3C_142_gat) );
BUFX20 U_g247 (.A(GS3_117_gat), .Y(GY3D_143_gat) );
BUFX20 U_g248 (.A(GS3_117_gat), .Y(GY3I_144_gat) );
BUFX20 U_g249 (.A(GS3_117_gat), .Y(GY3K_145_gat) );
BUFX20 U_g250 (.A(GS2_118_gat), .Y(GY2A_146_gat) );
BUFX20 U_g251 (.A(GS2_118_gat), .Y(GY2C_147_gat) );
BUFX20 U_g252 (.A(GS2_118_gat), .Y(GY2D_148_gat) );
BUFX20 U_g253 (.A(GS2_118_gat), .Y(GY2J_149_gat) );
BUFX20 U_g254 (.A(GS2_118_gat), .Y(GY2L_150_gat) );
BUFX20 U_g255 (.A(GS1_119_gat), .Y(GY1A_151_gat) );
BUFX20 U_g256 (.A(GS1_119_gat), .Y(GY1B_152_gat) );
BUFX20 U_g257 (.A(GS1_119_gat), .Y(GY1D_153_gat) );
BUFX20 U_g258 (.A(GS1_119_gat), .Y(GY1I_154_gat) );
BUFX20 U_g259 (.A(GS1_119_gat), .Y(GY1J_155_gat) );
BUFX20 U_g260 (.A(GS0_120_gat), .Y(GY0A_156_gat) );
BUFX20 U_g261 (.A(GS0_120_gat), .Y(GY0B_157_gat) );
BUFX20 U_g262 (.A(GS0_120_gat), .Y(GY0C_158_gat) );
BUFX20 U_g263 (.A(GS0_120_gat), .Y(GY0K_159_gat) );
BUFX20 U_g264 (.A(GS0_120_gat), .Y(GY0L_160_gat) );
AND4XL U_g265 (.A(GS7_113_gat), .B(GY6A_126_gat), .C(GY5A_131_gat), .D(GY4A_136_gat), .Y(GT4_161_gat) );
AND4XL U_g266 (.A(GY7B_121_gat), .B(GS6_114_gat), .C(GY5B_132_gat), .D(GY4B_137_gat), .Y(GT5_162_gat) );
AND4XL U_g267 (.A(GY7C_122_gat), .B(GY6C_127_gat), .C(GS5_115_gat), .D(GY4C_138_gat), .Y(GT6_163_gat) );
AND4XL U_g268 (.A(GY7D_123_gat), .B(GY6D_128_gat), .C(GY5D_133_gat), .D(GS4_116_gat), .Y(GT7_164_gat) );
AND4XL U_g269 (.A(GS3_117_gat), .B(GY2A_146_gat), .C(GY1A_151_gat), .D(GY0A_156_gat), .Y(GT0_165_gat) );
AND4XL U_g270 (.A(GY3B_141_gat), .B(GS2_118_gat), .C(GY1B_152_gat), .D(GY0B_157_gat), .Y(GT1_166_gat) );
AND4XL U_g271 (.A(GY3C_142_gat), .B(GY2C_147_gat), .C(GS1_119_gat), .D(GY0C_158_gat), .Y(GT2_167_gat) );
AND4XL U_g272 (.A(GY3D_143_gat), .B(GY2D_148_gat), .C(GY1D_153_gat), .D(GS0_120_gat), .Y(GT3_168_gat) );
AND4XL U_g273 (.A(GT7_164_ngat), .B(GT6_163_ngat), .C(GT5_162_ngat), .D(GT4_161_ngat), .Y(GU1_169_gat) );
AND4XL U_g274 (.A(GT3_168_ngat), .B(GT2_167_ngat), .C(GT1_166_ngat), .D(GT0_165_ngat), .Y(GU0_170_gat) );
AND5XL U_g275 (.A(GU0_170_gat), .B(GS7_113_gat), .C(GY6J_129_gat), .D(GY5J_135_gat), .E(GS4_116_gat), .Y(GWB_171_gat) );
AND5XL U_g276 (.A(GU0_170_gat), .B(GS7_113_gat), .C(GY6L_130_gat), .D(GS5_115_gat), .E(GY4L_140_gat), .Y(GWD_172_gat) );
AND5XL U_g277 (.A(GU0_170_gat), .B(GY7I_124_gat), .C(GS6_114_gat), .D(GY5I_134_gat), .E(GS4_116_gat), .Y(GWA_173_gat) );
AND5XL U_g278 (.A(GU0_170_gat), .B(GY7K_125_gat), .C(GS6_114_gat), .D(GS5_115_gat), .E(GY4K_139_gat), .Y(GWC_174_gat) );
AND5XL U_g279 (.A(GU1_169_gat), .B(GS3_117_gat), .C(GY2J_149_gat), .D(GY1J_155_gat), .E(GS0_120_gat), .Y(GWF_175_gat) );
AND5XL U_g280 (.A(GU1_169_gat), .B(GS3_117_gat), .C(GY2L_150_gat), .D(GS1_119_gat), .E(GY0L_160_gat), .Y(GWH_176_gat) );
AND5XL U_g281 (.A(GU1_169_gat), .B(GY3I_144_gat), .C(GS2_118_gat), .D(GY1I_154_gat), .E(GS0_120_gat), .Y(GWE_177_gat) );
AND5XL U_g282 (.A(GU1_169_gat), .B(GY3K_145_gat), .C(GS2_118_gat), .D(GS1_119_gat), .E(GY0K_159_gat), .Y(GWG_178_gat) );
AND2XL U_g283 (.A(GWE_177_gat), .B(GS7_113_gat), .Y(GE19_179_gat) );
AND2XL U_g284 (.A(GWF_175_gat), .B(GS7_113_gat), .Y(GE23_180_gat) );
AND2XL U_g285 (.A(GWG_178_gat), .B(GS7_113_gat), .Y(GE27_181_gat) );
AND2XL U_g286 (.A(GWH_176_gat), .B(GS7_113_gat), .Y(GE31_182_gat) );
AND2XL U_g287 (.A(GWE_177_gat), .B(GS6_114_gat), .Y(GE18_183_gat) );
AND2XL U_g288 (.A(GWF_175_gat), .B(GS6_114_gat), .Y(GE22_184_gat) );
AND2XL U_g289 (.A(GWG_178_gat), .B(GS6_114_gat), .Y(GE26_185_gat) );
AND2XL U_g290 (.A(GWH_176_gat), .B(GS6_114_gat), .Y(GE30_186_gat) );
AND2XL U_g291 (.A(GWE_177_gat), .B(GS5_115_gat), .Y(GE17_187_gat) );
AND2XL U_g292 (.A(GWF_175_gat), .B(GS5_115_gat), .Y(GE21_188_gat) );
AND2XL U_g293 (.A(GWG_178_gat), .B(GS5_115_gat), .Y(GE25_189_gat) );
AND2XL U_g294 (.A(GWH_176_gat), .B(GS5_115_gat), .Y(GE29_190_gat) );
AND2XL U_g295 (.A(GWE_177_gat), .B(GS4_116_gat), .Y(GE16_191_gat) );
AND2XL U_g296 (.A(GWF_175_gat), .B(GS4_116_gat), .Y(GE20_192_gat) );
AND2XL U_g297 (.A(GWG_178_gat), .B(GS4_116_gat), .Y(GE24_193_gat) );
AND2XL U_g298 (.A(GWH_176_gat), .B(GS4_116_gat), .Y(GE28_194_gat) );
AND2XL U_g299 (.A(GWA_173_gat), .B(GS3_117_gat), .Y(GE3_195_gat) );
AND2XL U_g300 (.A(GWB_171_gat), .B(GS3_117_gat), .Y(GE7_196_gat) );
AND2XL U_g301 (.A(GWC_174_gat), .B(GS3_117_gat), .Y(GE11_197_gat) );
AND2XL U_g302 (.A(GWD_172_gat), .B(GS3_117_gat), .Y(GE15_198_gat) );
AND2XL U_g303 (.A(GWA_173_gat), .B(GS2_118_gat), .Y(GE2_199_gat) );
AND2XL U_g304 (.A(GWB_171_gat), .B(GS2_118_gat), .Y(GE6_200_gat) );
AND2XL U_g305 (.A(GWC_174_gat), .B(GS2_118_gat), .Y(GE10_201_gat) );
AND2XL U_g306 (.A(GWD_172_gat), .B(GS2_118_gat), .Y(GE14_202_gat) );
AND2XL U_g307 (.A(GWA_173_gat), .B(GS1_119_gat), .Y(GE1_203_gat) );
AND2XL U_g308 (.A(GWB_171_gat), .B(GS1_119_gat), .Y(GE5_204_gat) );
AND2XL U_g309 (.A(GWC_174_gat), .B(GS1_119_gat), .Y(GE9_205_gat) );
AND2XL U_g310 (.A(GWD_172_gat), .B(GS1_119_gat), .Y(GE13_206_gat) );
AND2XL U_g311 (.A(GWA_173_gat), .B(GS0_120_gat), .Y(GE0_207_gat) );
AND2XL U_g312 (.A(GWB_171_gat), .B(GS0_120_gat), .Y(GE4_208_gat) );
AND2XL U_g313 (.A(GWC_174_gat), .B(GS0_120_gat), .Y(GE8_209_gat) );
AND2XL U_g314 (.A(GWD_172_gat), .B(GS0_120_gat), .Y(GE12_210_gat) );
OR2XL U_g315 (.A(Ginternal__317gat), .B(Ginternal__316gat), .Y(GOD31_211_gat) );
AND2XL U_g316 (.A(GE31_182_gat), .B(GID31_31_ngat), .Y(Ginternal__316gat) );
AND2XL U_g317 (.A(GE31_182_ngat), .B(GID31_31_gat), .Y(Ginternal__317gat) );
OR2XL U_g318 (.A(Ginternal__320gat), .B(Ginternal__319gat), .Y(GOD30_212_gat) );
AND2XL U_g319 (.A(GE30_186_gat), .B(GID30_30_ngat), .Y(Ginternal__319gat) );
AND2XL U_g320 (.A(GE30_186_ngat), .B(GID30_30_gat), .Y(Ginternal__320gat) );
OR2XL U_g321 (.A(Ginternal__323gat), .B(Ginternal__322gat), .Y(GOD29_213_gat) );
AND2XL U_g322 (.A(GE29_190_gat), .B(GID29_29_ngat), .Y(Ginternal__322gat) );
AND2XL U_g323 (.A(GE29_190_ngat), .B(GID29_29_gat), .Y(Ginternal__323gat) );
OR2XL U_g324 (.A(Ginternal__326gat), .B(Ginternal__325gat), .Y(GOD28_214_gat) );
AND2XL U_g325 (.A(GE28_194_gat), .B(GID28_28_ngat), .Y(Ginternal__325gat) );
AND2XL U_g326 (.A(GE28_194_ngat), .B(GID28_28_gat), .Y(Ginternal__326gat) );
OR2XL U_g327 (.A(Ginternal__329gat), .B(Ginternal__328gat), .Y(GOD27_215_gat) );
AND2XL U_g328 (.A(GE27_181_gat), .B(GID27_27_ngat), .Y(Ginternal__328gat) );
AND2XL U_g329 (.A(GE27_181_ngat), .B(GID27_27_gat), .Y(Ginternal__329gat) );
OR2XL U_g330 (.A(Ginternal__332gat), .B(Ginternal__331gat), .Y(GOD26_216_gat) );
AND2XL U_g331 (.A(GE26_185_gat), .B(GID26_26_ngat), .Y(Ginternal__331gat) );
AND2XL U_g332 (.A(GE26_185_ngat), .B(GID26_26_gat), .Y(Ginternal__332gat) );
OR2XL U_g333 (.A(Ginternal__335gat), .B(Ginternal__334gat), .Y(GOD25_217_gat) );
AND2XL U_g334 (.A(GE25_189_gat), .B(GID25_25_ngat), .Y(Ginternal__334gat) );
AND2XL U_g335 (.A(GE25_189_ngat), .B(GID25_25_gat), .Y(Ginternal__335gat) );
OR2XL U_g336 (.A(Ginternal__338gat), .B(Ginternal__337gat), .Y(GOD24_218_gat) );
AND2XL U_g337 (.A(GE24_193_gat), .B(GID24_24_ngat), .Y(Ginternal__337gat) );
AND2XL U_g338 (.A(GE24_193_ngat), .B(GID24_24_gat), .Y(Ginternal__338gat) );
OR2XL U_g339 (.A(Ginternal__341gat), .B(Ginternal__340gat), .Y(GOD23_219_gat) );
AND2XL U_g340 (.A(GE23_180_gat), .B(GID23_23_ngat), .Y(Ginternal__340gat) );
AND2XL U_g341 (.A(GE23_180_ngat), .B(GID23_23_gat), .Y(Ginternal__341gat) );
OR2XL U_g342 (.A(Ginternal__344gat), .B(Ginternal__343gat), .Y(GOD22_220_gat) );
AND2XL U_g343 (.A(GE22_184_gat), .B(GID22_22_ngat), .Y(Ginternal__343gat) );
AND2XL U_g344 (.A(GE22_184_ngat), .B(GID22_22_gat), .Y(Ginternal__344gat) );
OR2XL U_g345 (.A(Ginternal__347gat), .B(Ginternal__346gat), .Y(GOD21_221_gat) );
AND2XL U_g346 (.A(GE21_188_gat), .B(GID21_21_ngat), .Y(Ginternal__346gat) );
AND2XL U_g347 (.A(GE21_188_ngat), .B(GID21_21_gat), .Y(Ginternal__347gat) );
OR2XL U_g348 (.A(Ginternal__350gat), .B(Ginternal__349gat), .Y(GOD20_222_gat) );
AND2XL U_g349 (.A(GE20_192_gat), .B(GID20_20_ngat), .Y(Ginternal__349gat) );
AND2XL U_g350 (.A(GE20_192_ngat), .B(GID20_20_gat), .Y(Ginternal__350gat) );
OR2XL U_g351 (.A(Ginternal__353gat), .B(Ginternal__352gat), .Y(GOD19_223_gat) );
AND2XL U_g352 (.A(GE19_179_gat), .B(GID19_19_ngat), .Y(Ginternal__352gat) );
AND2XL U_g353 (.A(GE19_179_ngat), .B(GID19_19_gat), .Y(Ginternal__353gat) );
OR2XL U_g354 (.A(Ginternal__356gat), .B(Ginternal__355gat), .Y(GOD18_224_gat) );
AND2XL U_g355 (.A(GE18_183_gat), .B(GID18_18_ngat), .Y(Ginternal__355gat) );
AND2XL U_g356 (.A(GE18_183_ngat), .B(GID18_18_gat), .Y(Ginternal__356gat) );
OR2XL U_g357 (.A(Ginternal__359gat), .B(Ginternal__358gat), .Y(GOD17_225_gat) );
AND2XL U_g358 (.A(GE17_187_gat), .B(GID17_17_ngat), .Y(Ginternal__358gat) );
AND2XL U_g359 (.A(GE17_187_ngat), .B(GID17_17_gat), .Y(Ginternal__359gat) );
OR2XL U_g360 (.A(Ginternal__362gat), .B(Ginternal__361gat), .Y(GOD16_226_gat) );
AND2XL U_g361 (.A(GE16_191_gat), .B(GID16_16_ngat), .Y(Ginternal__361gat) );
AND2XL U_g362 (.A(GE16_191_ngat), .B(GID16_16_gat), .Y(Ginternal__362gat) );
OR2XL U_g363 (.A(Ginternal__365gat), .B(Ginternal__364gat), .Y(GOD15_227_gat) );
AND2XL U_g364 (.A(GE15_198_gat), .B(GID15_15_ngat), .Y(Ginternal__364gat) );
AND2XL U_g365 (.A(GE15_198_ngat), .B(GID15_15_gat), .Y(Ginternal__365gat) );
OR2XL U_g366 (.A(Ginternal__368gat), .B(Ginternal__367gat), .Y(GOD14_228_gat) );
AND2XL U_g367 (.A(GE14_202_gat), .B(GID14_14_ngat), .Y(Ginternal__367gat) );
AND2XL U_g368 (.A(GE14_202_ngat), .B(GID14_14_gat), .Y(Ginternal__368gat) );
OR2XL U_g369 (.A(Ginternal__371gat), .B(Ginternal__370gat), .Y(GOD13_229_gat) );
AND2XL U_g370 (.A(GE13_206_gat), .B(GID13_13_ngat), .Y(Ginternal__370gat) );
AND2XL U_g371 (.A(GE13_206_ngat), .B(GID13_13_gat), .Y(Ginternal__371gat) );
OR2XL U_g372 (.A(Ginternal__374gat), .B(Ginternal__373gat), .Y(GOD12_230_gat) );
AND2XL U_g373 (.A(GE12_210_gat), .B(GID12_12_ngat), .Y(Ginternal__373gat) );
AND2XL U_g374 (.A(GE12_210_ngat), .B(GID12_12_gat), .Y(Ginternal__374gat) );
OR2XL U_g375 (.A(Ginternal__377gat), .B(Ginternal__376gat), .Y(GOD11_231_gat) );
AND2XL U_g376 (.A(GE11_197_gat), .B(GID11_11_ngat), .Y(Ginternal__376gat) );
AND2XL U_g377 (.A(GE11_197_ngat), .B(GID11_11_gat), .Y(Ginternal__377gat) );
OR2XL U_g378 (.A(Ginternal__380gat), .B(Ginternal__379gat), .Y(GOD10_232_gat) );
AND2XL U_g379 (.A(GE10_201_gat), .B(GID10_10_ngat), .Y(Ginternal__379gat) );
AND2XL U_g380 (.A(GE10_201_ngat), .B(GID10_10_gat), .Y(Ginternal__380gat) );
OR2XL U_g381 (.A(Ginternal__383gat), .B(Ginternal__382gat), .Y(GOD9_233_gat) );
AND2XL U_g382 (.A(GE9_205_gat), .B(GID9_9_ngat), .Y(Ginternal__382gat) );
AND2XL U_g383 (.A(GE9_205_ngat), .B(GID9_9_gat), .Y(Ginternal__383gat) );
OR2XL U_g384 (.A(Ginternal__386gat), .B(Ginternal__385gat), .Y(GOD8_234_gat) );
AND2XL U_g385 (.A(GE8_209_gat), .B(GID8_8_ngat), .Y(Ginternal__385gat) );
AND2XL U_g386 (.A(GE8_209_ngat), .B(GID8_8_gat), .Y(Ginternal__386gat) );
OR2XL U_g387 (.A(Ginternal__389gat), .B(Ginternal__388gat), .Y(GOD7_235_gat) );
AND2XL U_g388 (.A(GE7_196_gat), .B(GID7_7_ngat), .Y(Ginternal__388gat) );
AND2XL U_g389 (.A(GE7_196_ngat), .B(GID7_7_gat), .Y(Ginternal__389gat) );
OR2XL U_g390 (.A(Ginternal__392gat), .B(Ginternal__391gat), .Y(GOD6_236_gat) );
AND2XL U_g391 (.A(GE6_200_gat), .B(GID6_6_ngat), .Y(Ginternal__391gat) );
AND2XL U_g392 (.A(GE6_200_ngat), .B(GID6_6_gat), .Y(Ginternal__392gat) );
OR2XL U_g393 (.A(Ginternal__395gat), .B(Ginternal__394gat), .Y(GOD5_237_gat) );
AND2XL U_g394 (.A(GE5_204_gat), .B(GID5_5_ngat), .Y(Ginternal__394gat) );
AND2XL U_g395 (.A(GE5_204_ngat), .B(GID5_5_gat), .Y(Ginternal__395gat) );
OR2XL U_g396 (.A(Ginternal__398gat), .B(Ginternal__397gat), .Y(GOD4_238_gat) );
AND2XL U_g397 (.A(GE4_208_gat), .B(GID4_4_ngat), .Y(Ginternal__397gat) );
AND2XL U_g398 (.A(GE4_208_ngat), .B(GID4_4_gat), .Y(Ginternal__398gat) );
OR2XL U_g399 (.A(Ginternal__401gat), .B(Ginternal__400gat), .Y(GOD3_239_gat) );
AND2XL U_g400 (.A(GE3_195_gat), .B(GID3_3_ngat), .Y(Ginternal__400gat) );
AND2XL U_g401 (.A(GE3_195_ngat), .B(GID3_3_gat), .Y(Ginternal__401gat) );
OR2XL U_g402 (.A(Ginternal__404gat), .B(Ginternal__403gat), .Y(GOD2_240_gat) );
AND2XL U_g403 (.A(GE2_199_gat), .B(GID2_2_ngat), .Y(Ginternal__403gat) );
AND2XL U_g404 (.A(GE2_199_ngat), .B(GID2_2_gat), .Y(Ginternal__404gat) );
OR2XL U_g405 (.A(Ginternal__407gat), .B(Ginternal__406gat), .Y(GOD1_241_gat) );
AND2XL U_g406 (.A(GE1_203_gat), .B(GID1_1_ngat), .Y(Ginternal__406gat) );
AND2XL U_g407 (.A(GE1_203_ngat), .B(GID1_1_gat), .Y(Ginternal__407gat) );
OR2XL U_g408 (.A(Ginternal__410gat), .B(Ginternal__409gat), .Y(GOD0_242_gat) );
AND2XL U_g409 (.A(GE0_207_gat), .B(GID0_0_ngat), .Y(Ginternal__409gat) );
AND2XL U_g410 (.A(GE0_207_ngat), .B(GID0_0_gat), .Y(Ginternal__410gat) );
INVXL U_g411 (.A(GID30_30_gat), .Y(GID30_30_ngat) );
INVXL U_g412 (.A(GID31_31_gat), .Y(GID31_31_ngat) );
INVXL U_g413 (.A(GID28_28_gat), .Y(GID28_28_ngat) );
INVXL U_g414 (.A(GID29_29_gat), .Y(GID29_29_ngat) );
INVXL U_g415 (.A(GID27_27_gat), .Y(GID27_27_ngat) );
INVXL U_g416 (.A(GID26_26_gat), .Y(GID26_26_ngat) );
INVXL U_g417 (.A(GID25_25_gat), .Y(GID25_25_ngat) );
INVXL U_g418 (.A(GID24_24_gat), .Y(GID24_24_ngat) );
INVXL U_g419 (.A(GID22_22_gat), .Y(GID22_22_ngat) );
INVXL U_g420 (.A(GID23_23_gat), .Y(GID23_23_ngat) );
INVXL U_g421 (.A(GID20_20_gat), .Y(GID20_20_ngat) );
INVXL U_g422 (.A(GID21_21_gat), .Y(GID21_21_ngat) );
INVXL U_g423 (.A(GID19_19_gat), .Y(GID19_19_ngat) );
INVXL U_g424 (.A(GID18_18_gat), .Y(GID18_18_ngat) );
INVXL U_g425 (.A(GID17_17_gat), .Y(GID17_17_ngat) );
INVXL U_g426 (.A(GID16_16_gat), .Y(GID16_16_ngat) );
INVXL U_g427 (.A(GID14_14_gat), .Y(GID14_14_ngat) );
INVXL U_g428 (.A(GID15_15_gat), .Y(GID15_15_ngat) );
INVXL U_g429 (.A(GID12_12_gat), .Y(GID12_12_ngat) );
INVXL U_g430 (.A(GID13_13_gat), .Y(GID13_13_ngat) );
INVXL U_g431 (.A(GID11_11_gat), .Y(GID11_11_ngat) );
INVXL U_g432 (.A(GID10_10_gat), .Y(GID10_10_ngat) );
INVXL U_g433 (.A(GID9_9_gat), .Y(GID9_9_ngat) );
INVXL U_g434 (.A(GID8_8_gat), .Y(GID8_8_ngat) );
INVXL U_g435 (.A(GID6_6_gat), .Y(GID6_6_ngat) );
INVXL U_g436 (.A(GID7_7_gat), .Y(GID7_7_ngat) );
INVXL U_g437 (.A(GID4_4_gat), .Y(GID4_4_ngat) );
INVXL U_g438 (.A(GID5_5_gat), .Y(GID5_5_ngat) );
INVXL U_g439 (.A(GID3_3_gat), .Y(GID3_3_ngat) );
INVXL U_g440 (.A(GID2_2_gat), .Y(GID2_2_ngat) );
INVXL U_g441 (.A(GID1_1_gat), .Y(GID1_1_ngat) );
INVXL U_g442 (.A(GID0_0_gat), .Y(GID0_0_ngat) );
INVXL U_g443 (.A(GXA14_50_gat), .Y(GXA14_50_ngat) );
INVXL U_g444 (.A(GXA15_49_gat), .Y(GXA15_49_ngat) );
INVXL U_g445 (.A(GXB7_59_gat), .Y(GXB7_59_ngat) );
INVXL U_g446 (.A(GXC7_51_gat), .Y(GXC7_51_ngat) );
INVXL U_g447 (.A(GXB6_60_gat), .Y(GXB6_60_ngat) );
INVXL U_g448 (.A(GXC6_52_gat), .Y(GXC6_52_ngat) );
INVXL U_g449 (.A(GXA12_56_gat), .Y(GXA12_56_ngat) );
INVXL U_g450 (.A(GXA13_53_gat), .Y(GXA13_53_ngat) );
INVXL U_g451 (.A(GXB5_62_gat), .Y(GXB5_62_ngat) );
INVXL U_g452 (.A(GXC5_54_gat), .Y(GXC5_54_ngat) );
INVXL U_g453 (.A(GXB4_63_gat), .Y(GXB4_63_ngat) );
INVXL U_g454 (.A(GXC4_55_gat), .Y(GXC4_55_ngat) );
INVXL U_g455 (.A(GXA10_58_gat), .Y(GXA10_58_ngat) );
INVXL U_g456 (.A(GXA11_57_gat), .Y(GXA11_57_ngat) );
INVXL U_g457 (.A(GXA8_64_gat), .Y(GXA8_64_ngat) );
INVXL U_g458 (.A(GXA9_61_gat), .Y(GXA9_61_ngat) );
INVXL U_g459 (.A(GXA6_66_gat), .Y(GXA6_66_ngat) );
INVXL U_g460 (.A(GXA7_65_gat), .Y(GXA7_65_ngat) );
INVXL U_g461 (.A(GXB3_75_gat), .Y(GXB3_75_ngat) );
INVXL U_g462 (.A(GXC3_67_gat), .Y(GXC3_67_ngat) );
INVXL U_g463 (.A(GXB2_76_gat), .Y(GXB2_76_ngat) );
INVXL U_g464 (.A(GXC2_68_gat), .Y(GXC2_68_ngat) );
INVXL U_g465 (.A(GXA4_72_gat), .Y(GXA4_72_ngat) );
INVXL U_g466 (.A(GXA5_69_gat), .Y(GXA5_69_ngat) );
INVXL U_g467 (.A(GXB1_78_gat), .Y(GXB1_78_ngat) );
INVXL U_g468 (.A(GXC1_70_gat), .Y(GXC1_70_ngat) );
INVXL U_g469 (.A(GXB0_79_gat), .Y(GXB0_79_ngat) );
INVXL U_g470 (.A(GXC0_71_gat), .Y(GXC0_71_ngat) );
INVXL U_g471 (.A(GXA2_74_gat), .Y(GXA2_74_ngat) );
INVXL U_g472 (.A(GXA3_73_gat), .Y(GXA3_73_ngat) );
INVXL U_g473 (.A(GXA0_80_gat), .Y(GXA0_80_ngat) );
INVXL U_g474 (.A(GXA1_77_gat), .Y(GXA1_77_ngat) );
INVXL U_g475 (.A(GF6_84_gat), .Y(GF6_84_ngat) );
INVXL U_g476 (.A(GF7_81_gat), .Y(GF7_81_ngat) );
INVXL U_g477 (.A(GF5_87_gat), .Y(GF5_87_ngat) );
INVXL U_g478 (.A(GF4_88_gat), .Y(GF4_88_ngat) );
INVXL U_g479 (.A(GF2_92_gat), .Y(GF2_92_ngat) );
INVXL U_g480 (.A(GF3_89_gat), .Y(GF3_89_ngat) );
INVXL U_g481 (.A(GF1_95_gat), .Y(GF1_95_ngat) );
INVXL U_g482 (.A(GF0_96_gat), .Y(GF0_96_ngat) );
INVXL U_g483 (.A(GH7_41_gat), .Y(GH7_41_ngat) );
INVXL U_g484 (.A(GG3_102_gat), .Y(GG3_102_ngat) );
INVXL U_g485 (.A(GH6_42_gat), .Y(GH6_42_ngat) );
INVXL U_g486 (.A(GG2_103_gat), .Y(GG2_103_ngat) );
INVXL U_g487 (.A(GH5_43_gat), .Y(GH5_43_ngat) );
INVXL U_g488 (.A(GG1_101_gat), .Y(GG1_101_ngat) );
INVXL U_g489 (.A(GH4_44_gat), .Y(GH4_44_ngat) );
INVXL U_g490 (.A(GG0_104_gat), .Y(GG0_104_ngat) );
INVXL U_g491 (.A(GH3_45_gat), .Y(GH3_45_ngat) );
INVXL U_g492 (.A(GG7_98_gat), .Y(GG7_98_ngat) );
INVXL U_g493 (.A(GH2_46_gat), .Y(GH2_46_ngat) );
INVXL U_g494 (.A(GG6_99_gat), .Y(GG6_99_ngat) );
INVXL U_g495 (.A(GH1_47_gat), .Y(GH1_47_ngat) );
INVXL U_g496 (.A(GG5_97_gat), .Y(GG5_97_ngat) );
INVXL U_g497 (.A(GH0_48_gat), .Y(GH0_48_ngat) );
INVXL U_g498 (.A(GG4_100_gat), .Y(GG4_100_ngat) );
INVXL U_g499 (.A(GXE7_82_gat), .Y(GXE7_82_ngat) );
INVXL U_g500 (.A(GXD7_105_gat), .Y(GXD7_105_ngat) );
INVXL U_g501 (.A(GXE6_83_gat), .Y(GXE6_83_ngat) );
INVXL U_g502 (.A(GXD6_106_gat), .Y(GXD6_106_ngat) );
INVXL U_g503 (.A(GXE5_85_gat), .Y(GXE5_85_ngat) );
INVXL U_g504 (.A(GXD5_107_gat), .Y(GXD5_107_ngat) );
INVXL U_g505 (.A(GXE4_86_gat), .Y(GXE4_86_ngat) );
INVXL U_g506 (.A(GXD4_108_gat), .Y(GXD4_108_ngat) );
INVXL U_g507 (.A(GXE3_90_gat), .Y(GXE3_90_ngat) );
INVXL U_g508 (.A(GXD3_109_gat), .Y(GXD3_109_ngat) );
INVXL U_g509 (.A(GXE2_91_gat), .Y(GXE2_91_ngat) );
INVXL U_g510 (.A(GXD2_110_gat), .Y(GXD2_110_ngat) );
INVXL U_g511 (.A(GXE1_93_gat), .Y(GXE1_93_ngat) );
INVXL U_g512 (.A(GXD1_111_gat), .Y(GXD1_111_ngat) );
INVXL U_g513 (.A(GXE0_94_gat), .Y(GXE0_94_ngat) );
INVXL U_g514 (.A(GXD0_112_gat), .Y(GXD0_112_ngat) );
INVXL U_g515 (.A(GT4_161_gat), .Y(GT4_161_ngat) );
INVXL U_g516 (.A(GT5_162_gat), .Y(GT5_162_ngat) );
INVXL U_g517 (.A(GT6_163_gat), .Y(GT6_163_ngat) );
INVXL U_g518 (.A(GT7_164_gat), .Y(GT7_164_ngat) );
INVXL U_g519 (.A(GT0_165_gat), .Y(GT0_165_ngat) );
INVXL U_g520 (.A(GT1_166_gat), .Y(GT1_166_ngat) );
INVXL U_g521 (.A(GT2_167_gat), .Y(GT2_167_ngat) );
INVXL U_g522 (.A(GT3_168_gat), .Y(GT3_168_ngat) );
INVXL U_g523 (.A(GE31_182_gat), .Y(GE31_182_ngat) );
INVXL U_g524 (.A(GE30_186_gat), .Y(GE30_186_ngat) );
INVXL U_g525 (.A(GE29_190_gat), .Y(GE29_190_ngat) );
INVXL U_g526 (.A(GE28_194_gat), .Y(GE28_194_ngat) );
INVXL U_g527 (.A(GE27_181_gat), .Y(GE27_181_ngat) );
INVXL U_g528 (.A(GE26_185_gat), .Y(GE26_185_ngat) );
INVXL U_g529 (.A(GE25_189_gat), .Y(GE25_189_ngat) );
INVXL U_g530 (.A(GE24_193_gat), .Y(GE24_193_ngat) );
INVXL U_g531 (.A(GE23_180_gat), .Y(GE23_180_ngat) );
INVXL U_g532 (.A(GE22_184_gat), .Y(GE22_184_ngat) );
INVXL U_g533 (.A(GE21_188_gat), .Y(GE21_188_ngat) );
INVXL U_g534 (.A(GE20_192_gat), .Y(GE20_192_ngat) );
INVXL U_g535 (.A(GE19_179_gat), .Y(GE19_179_ngat) );
INVXL U_g536 (.A(GE18_183_gat), .Y(GE18_183_ngat) );
INVXL U_g537 (.A(GE17_187_gat), .Y(GE17_187_ngat) );
INVXL U_g538 (.A(GE16_191_gat), .Y(GE16_191_ngat) );
INVXL U_g539 (.A(GE15_198_gat), .Y(GE15_198_ngat) );
INVXL U_g540 (.A(GE14_202_gat), .Y(GE14_202_ngat) );
INVXL U_g541 (.A(GE13_206_gat), .Y(GE13_206_ngat) );
INVXL U_g542 (.A(GE12_210_gat), .Y(GE12_210_ngat) );
INVXL U_g543 (.A(GE11_197_gat), .Y(GE11_197_ngat) );
INVXL U_g544 (.A(GE10_201_gat), .Y(GE10_201_ngat) );
INVXL U_g545 (.A(GE9_205_gat), .Y(GE9_205_ngat) );
INVXL U_g546 (.A(GE8_209_gat), .Y(GE8_209_ngat) );
INVXL U_g547 (.A(GE7_196_gat), .Y(GE7_196_ngat) );
INVXL U_g548 (.A(GE6_200_gat), .Y(GE6_200_ngat) );
INVXL U_g549 (.A(GE5_204_gat), .Y(GE5_204_ngat) );
INVXL U_g550 (.A(GE4_208_gat), .Y(GE4_208_ngat) );
INVXL U_g551 (.A(GE3_195_gat), .Y(GE3_195_ngat) );
INVXL U_g552 (.A(GE2_199_gat), .Y(GE2_199_ngat) );
INVXL U_g553 (.A(GE1_203_gat), .Y(GE1_203_ngat) );
INVXL U_g554 (.A(GE0_207_gat), .Y(GE0_207_ngat) );

endmodule
