module C7552 ( G1_0_gat, G5_1_gat, G9_2_gat, G12_3_gat, G15_4_gat, G18_5_gat, G23_6_gat, G26_7_gat, G29_8_gat, G32_9_gat, G35_10_gat, G38_11_gat, G41_12_gat, G44_13_gat, G47_14_gat, G50_15_gat, G53_16_gat, G54_17_gat, G55_18_gat, G56_19_gat, G57_20_gat, G58_21_gat, G59_22_gat, G60_23_gat, G61_24_gat, G62_25_gat, G63_26_gat, G64_27_gat, G65_28_gat, G66_29_gat, G69_30_gat, G70_31_gat, G73_32_gat, G74_33_gat, G75_34_gat, G76_35_gat, G77_36_gat, G78_37_gat, G79_38_gat, G80_39_gat, G81_40_gat, G82_41_gat, G83_42_gat, G84_43_gat, G85_44_gat, G86_45_gat, G87_46_gat, G88_47_gat, G89_48_gat, G94_49_gat, G97_50_gat, G100_51_gat, G103_52_gat, G106_53_gat, G109_54_gat, G110_55_gat, G111_56_gat, G112_57_gat, G113_58_gat, G114_59_gat, G115_60_gat, G118_61_gat, G121_62_gat, G124_63_gat, G127_64_gat, G130_65_gat, G133_66_gat, G134_67_gat, G135_68_gat, G138_69_gat, G141_70_gat, G144_71_gat, G147_72_gat, G150_73_gat, G151_74_gat, G152_75_gat, G153_76_gat, G154_77_gat, G155_78_gat, G156_79_gat, G157_80_gat, G158_81_gat, G159_82_gat, G160_83_gat, G161_84_gat, G162_85_gat, G163_86_gat, G164_87_gat, G165_88_gat, G166_89_gat, G167_90_gat, G168_91_gat, G169_92_gat, G170_93_gat, G171_94_gat, G172_95_gat, G173_96_gat, G174_97_gat, G175_98_gat, G176_99_gat, G177_100_gat, G178_101_gat, G179_102_gat, G180_103_gat, G181_104_gat, G182_105_gat, G183_106_gat, G184_107_gat, G185_108_gat, G186_109_gat, G187_110_gat, G188_111_gat, G189_112_gat, G190_113_gat, G191_114_gat, G192_115_gat, G193_116_gat, G194_117_gat, G195_118_gat, G196_119_gat, G197_120_gat, G198_121_gat, G199_122_gat, G200_123_gat, G201_124_gat, G202_125_gat, G203_126_gat, G204_127_gat, G205_128_gat, G206_129_gat, G207_130_gat, G208_131_gat, G209_132_gat, G210_133_gat, G211_134_gat, G212_135_gat, G213_136_gat, G214_137_gat, G215_138_gat, G216_139_gat, G217_140_gat, G218_141_gat, G219_142_gat, G220_143_gat, G221_144_gat, G222_145_gat, G223_146_gat, G224_147_gat, G225_148_gat, G226_149_gat, G227_150_gat, G228_151_gat, G229_152_gat, G230_153_gat, G231_154_gat, G232_155_gat, G233_156_gat, G234_157_gat, G235_158_gat, G236_159_gat, G237_160_gat, G238_161_gat, G239_162_gat, G240_163_gat, GIN_339_164_gat, G1197_165_gat, G1455_166_gat, G1459_167_gat, G1462_168_gat, G1469_169_gat, G1480_170_gat, G1486_171_gat, G1492_172_gat, G1496_173_gat, G2204_174_gat, G2208_175_gat, G2211_176_gat, G2218_177_gat, G2224_178_gat, G2230_179_gat, G2236_180_gat, G2239_181_gat, G2247_182_gat, G2253_183_gat, G2256_184_gat, G3698_185_gat, G3701_186_gat, G3705_187_gat, G3711_188_gat, G3717_189_gat, G3723_190_gat, G3729_191_gat, G3737_192_gat, G3743_193_gat, G3749_194_gat, G4393_195_gat, G4394_196_gat, G4400_197_gat, G4405_198_gat, G4410_199_gat, G4415_200_gat, G4420_201_gat, G4427_202_gat, G4432_203_gat, G4437_204_gat, G4526_205_gat, G4528_206_gat, G339_164_gat, G2_313_gat, G3_312_gat, G450_288_gat, G448_284_gat, G444_282_gat, G442_280_gat, G440_277_gat, G438_274_gat, G496_271_gat, G494_267_gat, G492_265_gat, G490_263_gat, G488_260_gat, G486_258_gat, G484_256_gat, G482_253_gat, G480_250_gat, G560_248_gat, G542_246_gat, G558_244_gat, G556_242_gat, G554_240_gat, G552_238_gat, G550_236_gat, G548_234_gat, G546_232_gat, G544_230_gat, G540_227_gat, G538_224_gat, G536_222_gat, G534_220_gat, G532_218_gat, G530_216_gat, G528_214_gat, G526_212_gat, G524_210_gat, G279_304_gat, G436_286_gat, G478_269_gat, G522_226_gat, G402_395_gat, G404_390_gat, G406_388_gat, G408_385_gat, G410_387_gat, G432_428_gat, G446_393_gat, G284_384_gat, G286_419_gat, G289_383_gat, G292_392_gat, G341_420_gat, G281_547_gat, G453_596_gat, G278_536_gat, G373_2994_gat, G246_3110_gat, G258_3122_gat, G264_3121_gat, G270_3109_gat, G388_3093_gat, G391_3094_gat, G394_3095_gat, G397_3097_gat, G376_3206_gat, G379_3207_gat, G382_3148_gat, G385_3151_gat, G412_3369_gat, G414_3338_gat, G416_3368_gat, G249_3418_gat, G295_3352_gat, G324_3363_gat, G252_3450_gat, G276_3401_gat, G310_3393_gat, G313_3396_gat, G316_3397_gat, G319_3398_gat, G327_3408_gat, G330_3411_gat, G333_3416_gat, G336_3412_gat, G418_3449_gat, G273_3402_gat, G298_3387_gat, G301_3388_gat, G304_3390_gat, G307_3389_gat, G344_3382_gat, G422_3451_gat, G469_3452_gat, G419_3444_gat, G471_3445_gat, G359_3426_gat, G362_3429_gat, G365_3430_gat, G368_3431_gat, G347_3420_gat, G350_3421_gat, G353_3425_gat, G356_3424_gat, G321_3715_gat, G338_3716_gat, G370_3718_gat, G399_3717_gat);

input G1_0_gat;
input G5_1_gat;
input G9_2_gat;
input G12_3_gat;
input G15_4_gat;
input G18_5_gat;
input G23_6_gat;
input G26_7_gat;
input G29_8_gat;
input G32_9_gat;
input G35_10_gat;
input G38_11_gat;
input G41_12_gat;
input G44_13_gat;
input G47_14_gat;
input G50_15_gat;
input G53_16_gat;
input G54_17_gat;
input G55_18_gat;
input G56_19_gat;
input G57_20_gat;
input G58_21_gat;
input G59_22_gat;
input G60_23_gat;
input G61_24_gat;
input G62_25_gat;
input G63_26_gat;
input G64_27_gat;
input G65_28_gat;
input G66_29_gat;
input G69_30_gat;
input G70_31_gat;
input G73_32_gat;
input G74_33_gat;
input G75_34_gat;
input G76_35_gat;
input G77_36_gat;
input G78_37_gat;
input G79_38_gat;
input G80_39_gat;
input G81_40_gat;
input G82_41_gat;
input G83_42_gat;
input G84_43_gat;
input G85_44_gat;
input G86_45_gat;
input G87_46_gat;
input G88_47_gat;
input G89_48_gat;
input G94_49_gat;
input G97_50_gat;
input G100_51_gat;
input G103_52_gat;
input G106_53_gat;
input G109_54_gat;
input G110_55_gat;
input G111_56_gat;
input G112_57_gat;
input G113_58_gat;
input G114_59_gat;
input G115_60_gat;
input G118_61_gat;
input G121_62_gat;
input G124_63_gat;
input G127_64_gat;
input G130_65_gat;
input G133_66_gat;
input G134_67_gat;
input G135_68_gat;
input G138_69_gat;
input G141_70_gat;
input G144_71_gat;
input G147_72_gat;
input G150_73_gat;
input G151_74_gat;
input G152_75_gat;
input G153_76_gat;
input G154_77_gat;
input G155_78_gat;
input G156_79_gat;
input G157_80_gat;
input G158_81_gat;
input G159_82_gat;
input G160_83_gat;
input G161_84_gat;
input G162_85_gat;
input G163_86_gat;
input G164_87_gat;
input G165_88_gat;
input G166_89_gat;
input G167_90_gat;
input G168_91_gat;
input G169_92_gat;
input G170_93_gat;
input G171_94_gat;
input G172_95_gat;
input G173_96_gat;
input G174_97_gat;
input G175_98_gat;
input G176_99_gat;
input G177_100_gat;
input G178_101_gat;
input G179_102_gat;
input G180_103_gat;
input G181_104_gat;
input G182_105_gat;
input G183_106_gat;
input G184_107_gat;
input G185_108_gat;
input G186_109_gat;
input G187_110_gat;
input G188_111_gat;
input G189_112_gat;
input G190_113_gat;
input G191_114_gat;
input G192_115_gat;
input G193_116_gat;
input G194_117_gat;
input G195_118_gat;
input G196_119_gat;
input G197_120_gat;
input G198_121_gat;
input G199_122_gat;
input G200_123_gat;
input G201_124_gat;
input G202_125_gat;
input G203_126_gat;
input G204_127_gat;
input G205_128_gat;
input G206_129_gat;
input G207_130_gat;
input G208_131_gat;
input G209_132_gat;
input G210_133_gat;
input G211_134_gat;
input G212_135_gat;
input G213_136_gat;
input G214_137_gat;
input G215_138_gat;
input G216_139_gat;
input G217_140_gat;
input G218_141_gat;
input G219_142_gat;
input G220_143_gat;
input G221_144_gat;
input G222_145_gat;
input G223_146_gat;
input G224_147_gat;
input G225_148_gat;
input G226_149_gat;
input G227_150_gat;
input G228_151_gat;
input G229_152_gat;
input G230_153_gat;
input G231_154_gat;
input G232_155_gat;
input G233_156_gat;
input G234_157_gat;
input G235_158_gat;
input G236_159_gat;
input G237_160_gat;
input G238_161_gat;
input G239_162_gat;
input G240_163_gat;
input GIN_339_164_gat;
input G1197_165_gat;
input G1455_166_gat;
input G1459_167_gat;
input G1462_168_gat;
input G1469_169_gat;
input G1480_170_gat;
input G1486_171_gat;
input G1492_172_gat;
input G1496_173_gat;
input G2204_174_gat;
input G2208_175_gat;
input G2211_176_gat;
input G2218_177_gat;
input G2224_178_gat;
input G2230_179_gat;
input G2236_180_gat;
input G2239_181_gat;
input G2247_182_gat;
input G2253_183_gat;
input G2256_184_gat;
input G3698_185_gat;
input G3701_186_gat;
input G3705_187_gat;
input G3711_188_gat;
input G3717_189_gat;
input G3723_190_gat;
input G3729_191_gat;
input G3737_192_gat;
input G3743_193_gat;
input G3749_194_gat;
input G4393_195_gat;
input G4394_196_gat;
input G4400_197_gat;
input G4405_198_gat;
input G4410_199_gat;
input G4415_200_gat;
input G4420_201_gat;
input G4427_202_gat;
input G4432_203_gat;
input G4437_204_gat;
input G4526_205_gat;
input G4528_206_gat;

output G339_164_gat;
output G2_313_gat;
output G3_312_gat;
output G450_288_gat;
output G448_284_gat;
output G444_282_gat;
output G442_280_gat;
output G440_277_gat;
output G438_274_gat;
output G496_271_gat;
output G494_267_gat;
output G492_265_gat;
output G490_263_gat;
output G488_260_gat;
output G486_258_gat;
output G484_256_gat;
output G482_253_gat;
output G480_250_gat;
output G560_248_gat;
output G542_246_gat;
output G558_244_gat;
output G556_242_gat;
output G554_240_gat;
output G552_238_gat;
output G550_236_gat;
output G548_234_gat;
output G546_232_gat;
output G544_230_gat;
output G540_227_gat;
output G538_224_gat;
output G536_222_gat;
output G534_220_gat;
output G532_218_gat;
output G530_216_gat;
output G528_214_gat;
output G526_212_gat;
output G524_210_gat;
output G279_304_gat;
output G436_286_gat;
output G478_269_gat;
output G522_226_gat;
output G402_395_gat;
output G404_390_gat;
output G406_388_gat;
output G408_385_gat;
output G410_387_gat;
output G432_428_gat;
output G446_393_gat;
output G284_384_gat;
output G286_419_gat;
output G289_383_gat;
output G292_392_gat;
output G341_420_gat;
output G281_547_gat;
output G453_596_gat;
output G278_536_gat;
output G373_2994_gat;
output G246_3110_gat;
output G258_3122_gat;
output G264_3121_gat;
output G270_3109_gat;
output G388_3093_gat;
output G391_3094_gat;
output G394_3095_gat;
output G397_3097_gat;
output G376_3206_gat;
output G379_3207_gat;
output G382_3148_gat;
output G385_3151_gat;
output G412_3369_gat;
output G414_3338_gat;
output G416_3368_gat;
output G249_3418_gat;
output G295_3352_gat;
output G324_3363_gat;
output G252_3450_gat;
output G276_3401_gat;
output G310_3393_gat;
output G313_3396_gat;
output G316_3397_gat;
output G319_3398_gat;
output G327_3408_gat;
output G330_3411_gat;
output G333_3416_gat;
output G336_3412_gat;
output G418_3449_gat;
output G273_3402_gat;
output G298_3387_gat;
output G301_3388_gat;
output G304_3390_gat;
output G307_3389_gat;
output G344_3382_gat;
output G422_3451_gat;
output G469_3452_gat;
output G419_3444_gat;
output G471_3445_gat;
output G359_3426_gat;
output G362_3429_gat;
output G365_3430_gat;
output G368_3431_gat;
output G347_3420_gat;
output G350_3421_gat;
output G353_3425_gat;
output G356_3424_gat;
output G321_3715_gat;
output G338_3716_gat;
output G370_3718_gat;
output G399_3717_gat;

INVXL U_g1 (.A(G15_4_gat), .Y(G279_304_gat) );
OR2XL U_g2 (.A(G401_310_ngat), .B(G400_297_ngat), .Y(G402_395_gat) );
INVXL U_g3 (.A(G2857_293_gat), .Y(G404_390_gat) );
INVXL U_g4 (.A(G4514_292_gat), .Y(G406_388_gat) );
INVXL U_g5 (.A(G4442_290_gat), .Y(G408_385_gat) );
INVXL U_g6 (.A(G1501_291_gat), .Y(G410_387_gat) );
OR2XL U_g7 (.A(G574_308_ngat), .B(G1197_165_ngat), .Y(G284_384_gat) );
INVXL U_g8 (.A(G1205_305_gat), .Y(G286_419_gat) );
OR2XL U_g9 (.A(G574_308_ngat), .B(G1197_165_ngat), .Y(G289_383_gat) );
OR2XL U_g10 (.A(G575_309_ngat), .B(G1184_294_ngat), .Y(G292_392_gat) );
INVXL U_g11 (.A(G1205_305_gat), .Y(G341_420_gat) );
INVXL U_g12 (.A(G280_391_gat), .Y(G281_547_gat) );
AND2XL U_g13 (.A(G453_596_gat), .B(G163_86_gat), .Y(G278_536_gat) );
OR2XL U_g14 (.A(G372_2890_ngat), .B(G371_2754_ngat), .Y(G373_2994_gat) );
OR5XL U_g15 (.A(G245_2897_gat), .B(G244_3033_gat), .C(G243_3032_gat), .D(G242_2955_gat), .E(G241_2837_gat), .Y(G246_3110_gat) );
OR5XL U_g16 (.A(G257_2860_gat), .B(G256_2991_gat), .C(G255_2990_gat), .D(G254_2888_gat), .E(G3259_2874_gat), .Y(G258_3122_gat) );
OR5XL U_g17 (.A(G263_2858_gat), .B(G262_2993_gat), .C(G261_2992_gat), .D(G260_2889_gat), .E(G3259_2874_gat), .Y(G264_3121_gat) );
OR5XL U_g18 (.A(G269_2896_gat), .B(G268_3028_gat), .C(G267_3027_gat), .D(G266_2956_gat), .E(G265_2835_gat), .Y(G270_3109_gat) );
OR2XL U_g19 (.A(G387_2931_ngat), .B(G386_3020_ngat), .Y(G388_3093_gat) );
OR2XL U_g20 (.A(G390_2934_ngat), .B(G389_3021_ngat), .Y(G391_3094_gat) );
OR2XL U_g21 (.A(G393_2937_ngat), .B(G392_3022_ngat), .Y(G394_3095_gat) );
OR2XL U_g22 (.A(G396_2941_ngat), .B(G395_3023_ngat), .Y(G397_3097_gat) );
OR2XL U_g23 (.A(G375_3090_gat), .B(G374_3152_gat), .Y(G376_3206_gat) );
OR2XL U_g24 (.A(G378_3091_gat), .B(G377_3153_gat), .Y(G379_3207_gat) );
OR2XL U_g25 (.A(G381_3092_gat), .B(G380_3086_gat), .Y(G382_3148_gat) );
OR2XL U_g26 (.A(G384_3016_gat), .B(G383_3089_gat), .Y(G385_3151_gat) );
INVXL U_g27 (.A(G4443_3309_gat), .Y(G412_3369_gat) );
INVXL U_g28 (.A(G4524_3265_gat), .Y(G414_3338_gat) );
INVXL U_g29 (.A(G2868_3308_gat), .Y(G416_3368_gat) );
OR2XL U_g30 (.A(G248_3306_gat), .B(G247_3310_gat), .Y(G249_3418_gat) );
OR2XL U_g31 (.A(G294_3223_ngat), .B(G293_3285_ngat), .Y(G295_3352_gat) );
OR2XL U_g32 (.A(G323_3238_ngat), .B(G322_3302_ngat), .Y(G324_3363_gat) );
OR2XL U_g33 (.A(G251_3365_gat), .B(G250_3417_gat), .Y(G252_3450_gat) );
OR2XL U_g34 (.A(G275_3286_gat), .B(G274_3353_gat), .Y(G276_3401_gat) );
OR2XL U_g35 (.A(G309_3275_ngat), .B(G308_3346_ngat), .Y(G310_3393_gat) );
OR2XL U_g36 (.A(G312_3279_ngat), .B(G311_3349_ngat), .Y(G313_3396_gat) );
OR2XL U_g37 (.A(G315_3281_ngat), .B(G314_3350_ngat), .Y(G316_3397_gat) );
OR2XL U_g38 (.A(G318_3283_ngat), .B(G317_3351_ngat), .Y(G319_3398_gat) );
OR2XL U_g39 (.A(G326_3294_ngat), .B(G325_3358_ngat), .Y(G327_3408_gat) );
OR2XL U_g40 (.A(G329_3298_ngat), .B(G328_3361_ngat), .Y(G330_3411_gat) );
OR2XL U_g41 (.A(G332_3304_ngat), .B(G331_3364_ngat), .Y(G333_3416_gat) );
OR2XL U_g42 (.A(G335_3300_ngat), .B(G334_3362_ngat), .Y(G336_3412_gat) );
INVXL U_g43 (.A(G417_3415_gat), .Y(G418_3449_gat) );
OR2XL U_g44 (.A(G272_3287_gat), .B(G271_3354_gat), .Y(G273_3402_gat) );
OR2XL U_g45 (.A(G297_3266_gat), .B(G296_3340_gat), .Y(G298_3387_gat) );
OR2XL U_g46 (.A(G300_3267_gat), .B(G299_3341_gat), .Y(G301_3388_gat) );
OR2XL U_g47 (.A(G303_3271_gat), .B(G302_3342_gat), .Y(G304_3390_gat) );
OR2XL U_g48 (.A(G306_3270_gat), .B(G305_3343_gat), .Y(G307_3389_gat) );
OR2XL U_g49 (.A(G343_3258_ngat), .B(G342_3330_ngat), .Y(G344_3382_gat) );
OR2XL U_g50 (.A(G358_3320_ngat), .B(G357_3376_ngat), .Y(G359_3426_gat) );
OR2XL U_g51 (.A(G361_3324_ngat), .B(G360_3379_ngat), .Y(G362_3429_gat) );
OR2XL U_g52 (.A(G364_3326_ngat), .B(G363_3380_ngat), .Y(G365_3430_gat) );
OR2XL U_g53 (.A(G367_3328_ngat), .B(G366_3381_ngat), .Y(G368_3431_gat) );
OR2XL U_g54 (.A(G346_3311_gat), .B(G345_3370_gat), .Y(G347_3420_gat) );
OR2XL U_g55 (.A(G349_3314_gat), .B(G348_3371_gat), .Y(G350_3421_gat) );
OR2XL U_g56 (.A(G352_3318_gat), .B(G351_3372_gat), .Y(G353_3425_gat) );
OR2XL U_g57 (.A(G355_3317_gat), .B(G354_3375_gat), .Y(G356_3424_gat) );
INVXL U_g58 (.A(G320_3711_gat), .Y(G321_3715_gat) );
INVXL U_g59 (.A(G337_3712_gat), .Y(G338_3716_gat) );
INVXL U_g60 (.A(G369_3714_gat), .Y(G370_3718_gat) );
INVXL U_g61 (.A(G398_3713_gat), .Y(G399_3717_gat) );
BUFX20 U_g62 (.A(G4526_205_gat), .Y(G4833_207_gat) );
BUFX20 U_g63 (.A(G4526_205_gat), .Y(G2828_208_gat) );
INVXL U_g64 (.A(G4437_204_gat), .Y(G4439_209_gat) );
INVXL U_g65 (.A(G4432_203_gat), .Y(G4434_211_gat) );
INVXL U_g66 (.A(G4427_202_gat), .Y(G4429_213_gat) );
INVXL U_g67 (.A(G4420_201_gat), .Y(G4422_215_gat) );
INVXL U_g68 (.A(G4415_200_gat), .Y(G4417_217_gat) );
INVXL U_g69 (.A(G4410_199_gat), .Y(G4412_219_gat) );
INVXL U_g70 (.A(G4405_198_gat), .Y(G4407_221_gat) );
INVXL U_g71 (.A(G4400_197_gat), .Y(G4402_223_gat) );
INVXL U_g72 (.A(G4394_196_gat), .Y(G4396_225_gat) );
INVXL U_g73 (.A(G4393_195_gat), .Y(G4121_228_gat) );
INVXL U_g74 (.A(G3749_194_gat), .Y(G3751_229_gat) );
INVXL U_g75 (.A(G3743_193_gat), .Y(G3745_231_gat) );
INVXL U_g76 (.A(G3737_192_gat), .Y(G3739_233_gat) );
INVXL U_g77 (.A(G3729_191_gat), .Y(G3731_235_gat) );
INVXL U_g78 (.A(G3723_190_gat), .Y(G3725_237_gat) );
INVXL U_g79 (.A(G3717_189_gat), .Y(G3719_239_gat) );
INVXL U_g80 (.A(G3711_188_gat), .Y(G3713_241_gat) );
INVXL U_g81 (.A(G3705_187_gat), .Y(G3707_243_gat) );
INVXL U_g82 (.A(G3701_186_gat), .Y(G3703_245_gat) );
INVXL U_g83 (.A(G3698_185_gat), .Y(G3700_247_gat) );
INVXL U_g84 (.A(G2256_184_gat), .Y(G2258_249_gat) );
INVXL U_g85 (.A(G2256_184_gat), .Y(G1192_251_gat) );
INVXL U_g86 (.A(G2253_183_gat), .Y(G2255_252_gat) );
INVXL U_g87 (.A(G2253_183_gat), .Y(G1186_254_gat) );
INVXL U_g88 (.A(G2247_182_gat), .Y(G2249_255_gat) );
INVXL U_g89 (.A(G2239_181_gat), .Y(G2241_257_gat) );
INVXL U_g90 (.A(G2236_180_gat), .Y(G2238_259_gat) );
INVXL U_g91 (.A(G2236_180_gat), .Y(G1178_261_gat) );
INVXL U_g92 (.A(G2230_179_gat), .Y(G2232_262_gat) );
INVXL U_g93 (.A(G2224_178_gat), .Y(G2226_264_gat) );
INVXL U_g94 (.A(G2218_177_gat), .Y(G2220_266_gat) );
INVXL U_g95 (.A(G2211_176_gat), .Y(G2213_268_gat) );
INVXL U_g96 (.A(G2208_175_gat), .Y(G2210_270_gat) );
INVXL U_g97 (.A(G2204_174_gat), .Y(G2207_272_gat) );
INVXL U_g98 (.A(G1496_173_gat), .Y(G1499_273_gat) );
OR2XL U_g99 (.A(G1496_173_ngat), .B(G4528_206_ngat), .Y(G1541_275_gat) );
INVXL U_g100 (.A(G1492_172_gat), .Y(G1495_276_gat) );
AND2XL U_g101 (.A(G1492_172_gat), .B(G4528_206_gat), .Y(G1518_278_gat) );
INVXL U_g102 (.A(G1486_171_gat), .Y(G1488_279_gat) );
INVXL U_g103 (.A(G1480_170_gat), .Y(G1482_281_gat) );
INVXL U_g104 (.A(G1469_169_gat), .Y(G1471_283_gat) );
INVXL U_g105 (.A(G1462_168_gat), .Y(G1464_285_gat) );
INVXL U_g106 (.A(G1459_167_gat), .Y(G1461_287_gat) );
INVXL U_g107 (.A(G1455_166_gat), .Y(G1458_289_gat) );
AND4XL U_g108 (.A(G186_109_gat), .B(G185_108_gat), .C(G182_105_gat), .D(G183_106_gat), .Y(G4442_290_gat) );
AND4XL U_g109 (.A(G199_122_gat), .B(G188_111_gat), .C(G172_95_gat), .D(G162_85_gat), .Y(G1501_291_gat) );
AND4XL U_g110 (.A(G230_153_gat), .B(G218_141_gat), .C(G152_75_gat), .D(G210_133_gat), .Y(G4514_292_gat) );
AND4XL U_g111 (.A(G240_163_gat), .B(G228_151_gat), .C(G184_107_gat), .D(G150_73_gat), .Y(G2857_293_gat) );
AND2XL U_g112 (.A(G133_66_gat), .B(G134_67_gat), .Y(G1184_294_gat) );
BUFX20 U_g113 (.A(G106_53_gat), .Y(G446_393_gat) );
INVXL U_g114 (.A(G106_53_gat), .Y(G1500_296_gat) );
INVXL U_g115 (.A(G57_20_gat), .Y(G400_297_gat) );
BUFX20 U_g116 (.A(G38_11_gat), .Y(G1210_298_gat) );
BUFX20 U_g117 (.A(G38_11_gat), .Y(G1198_299_gat) );
BUFX20 U_g118 (.A(G18_5_gat), .Y(G1512_300_gat) );
BUFX20 U_g119 (.A(G18_5_gat), .Y(G1524_301_gat) );
INVXL U_g120 (.A(G18_5_gat), .Y(G1535_302_gat) );
BUFX20 U_g121 (.A(G18_5_gat), .Y(G1503_303_gat) );
BUFX20 U_g122 (.A(G15_4_gat), .Y(G1205_305_gat) );
OR2XL U_g123 (.A(G9_2_ngat), .B(G12_3_ngat), .Y(G1206_306_gat) );
OR2XL U_g124 (.A(G9_2_ngat), .B(G12_3_ngat), .Y(G1207_307_gat) );
INVXL U_g125 (.A(G5_1_gat), .Y(G574_308_gat) );
INVXL U_g126 (.A(G5_1_gat), .Y(G575_309_gat) );
INVXL U_g127 (.A(G5_1_gat), .Y(G401_310_gat) );
BUFX20 U_g128 (.A(G1_0_gat), .Y(G432_428_gat) );
OR2XL U_g129 (.A(G2207_272_ngat), .B(G4528_206_ngat), .Y(G2883_314_gat) );
AND2XL U_g130 (.A(G1458_289_gat), .B(G4528_206_gat), .Y(G2871_315_gat) );
INVXL U_g131 (.A(G4833_207_gat), .Y(G4839_316_gat) );
INVXL U_g132 (.A(G2828_208_gat), .Y(G2833_317_gat) );
BUFX20 U_g133 (.A(G4439_209_gat), .Y(G6853_318_gat) );
BUFX20 U_g134 (.A(G4439_209_gat), .Y(G6567_319_gat) );
BUFX20 U_g135 (.A(G4434_211_gat), .Y(G6575_320_gat) );
BUFX20 U_g136 (.A(G4434_211_gat), .Y(G6861_321_gat) );
BUFX20 U_g137 (.A(G4429_213_gat), .Y(G6583_322_gat) );
BUFX20 U_g138 (.A(G4429_213_gat), .Y(G6869_323_gat) );
BUFX20 U_g139 (.A(G4422_215_gat), .Y(G6909_324_gat) );
BUFX20 U_g140 (.A(G4422_215_gat), .Y(G6591_325_gat) );
BUFX20 U_g141 (.A(G4417_217_gat), .Y(G6877_326_gat) );
BUFX20 U_g142 (.A(G4417_217_gat), .Y(G6599_327_gat) );
BUFX20 U_g143 (.A(G4412_219_gat), .Y(G6607_328_gat) );
BUFX20 U_g144 (.A(G4412_219_gat), .Y(G6885_329_gat) );
BUFX20 U_g145 (.A(G4407_221_gat), .Y(G6893_330_gat) );
BUFX20 U_g146 (.A(G4407_221_gat), .Y(G6615_331_gat) );
BUFX20 U_g147 (.A(G4402_223_gat), .Y(G6901_332_gat) );
BUFX20 U_g148 (.A(G4402_223_gat), .Y(G6623_333_gat) );
BUFX20 U_g149 (.A(G4396_225_gat), .Y(G6631_334_gat) );
BUFX20 U_g150 (.A(G4396_225_gat), .Y(G6917_335_gat) );
BUFX20 U_g151 (.A(G3751_229_gat), .Y(G5985_336_gat) );
BUFX20 U_g152 (.A(G3751_229_gat), .Y(G5865_337_gat) );
BUFX20 U_g153 (.A(G3745_231_gat), .Y(G5873_338_gat) );
BUFX20 U_g154 (.A(G3745_231_gat), .Y(G5993_339_gat) );
BUFX20 U_g155 (.A(G3739_233_gat), .Y(G6001_340_gat) );
BUFX20 U_g156 (.A(G3739_233_gat), .Y(G5881_341_gat) );
BUFX20 U_g157 (.A(G3731_235_gat), .Y(G6041_342_gat) );
BUFX20 U_g158 (.A(G3731_235_gat), .Y(G5889_343_gat) );
BUFX20 U_g159 (.A(G3725_237_gat), .Y(G5897_344_gat) );
BUFX20 U_g160 (.A(G3725_237_gat), .Y(G6009_345_gat) );
BUFX20 U_g161 (.A(G3719_239_gat), .Y(G6017_346_gat) );
BUFX20 U_g162 (.A(G3719_239_gat), .Y(G5905_347_gat) );
BUFX20 U_g163 (.A(G3713_241_gat), .Y(G5913_348_gat) );
BUFX20 U_g164 (.A(G3713_241_gat), .Y(G6025_349_gat) );
BUFX20 U_g165 (.A(G3707_243_gat), .Y(G6033_350_gat) );
BUFX20 U_g166 (.A(G3707_243_gat), .Y(G5921_351_gat) );
BUFX20 U_g167 (.A(G1192_251_gat), .Y(G5393_352_gat) );
BUFX20 U_g168 (.A(G1192_251_gat), .Y(G5745_353_gat) );
BUFX20 U_g169 (.A(G1186_254_gat), .Y(G5753_354_gat) );
BUFX20 U_g170 (.A(G1186_254_gat), .Y(G5401_355_gat) );
BUFX20 U_g171 (.A(G2249_255_gat), .Y(G5409_356_gat) );
BUFX20 U_g172 (.A(G2249_255_gat), .Y(G5761_357_gat) );
BUFX20 U_g173 (.A(G2241_257_gat), .Y(G5769_358_gat) );
BUFX20 U_g174 (.A(G2241_257_gat), .Y(G5449_359_gat) );
BUFX20 U_g175 (.A(G1178_261_gat), .Y(G5417_360_gat) );
BUFX20 U_g176 (.A(G1178_261_gat), .Y(G5777_361_gat) );
BUFX20 U_g177 (.A(G2232_262_gat), .Y(G5785_362_gat) );
BUFX20 U_g178 (.A(G2232_262_gat), .Y(G5425_363_gat) );
BUFX20 U_g179 (.A(G2226_264_gat), .Y(G5433_364_gat) );
BUFX20 U_g180 (.A(G2226_264_gat), .Y(G5793_365_gat) );
BUFX20 U_g181 (.A(G2220_266_gat), .Y(G5801_366_gat) );
BUFX20 U_g182 (.A(G2220_266_gat), .Y(G5441_367_gat) );
BUFX20 U_g183 (.A(G2213_268_gat), .Y(G5457_368_gat) );
BUFX20 U_g184 (.A(G2213_268_gat), .Y(G5809_369_gat) );
AND2XL U_g185 (.A(G1198_299_gat), .B(G1541_275_gat), .Y(G777_370_gat) );
AND2XL U_g186 (.A(G1198_299_gat), .B(G1541_275_gat), .Y(G1115_371_gat) );
BUFX20 U_g187 (.A(G1541_275_gat), .Y(G5175_372_gat) );
BUFX20 U_g188 (.A(G1541_275_gat), .Y(G4873_373_gat) );
INVXL U_g189 (.A(G1518_278_gat), .Y(G1519_374_gat) );
BUFX20 U_g190 (.A(G1488_279_gat), .Y(G4881_375_gat) );
BUFX20 U_g191 (.A(G1488_279_gat), .Y(G5191_376_gat) );
BUFX20 U_g192 (.A(G1482_281_gat), .Y(G5199_377_gat) );
BUFX20 U_g193 (.A(G1482_281_gat), .Y(G4889_378_gat) );
BUFX20 U_g194 (.A(G1471_283_gat), .Y(G5215_379_gat) );
BUFX20 U_g195 (.A(G1471_283_gat), .Y(G4905_380_gat) );
BUFX20 U_g196 (.A(G1464_285_gat), .Y(G4921_381_gat) );
BUFX20 U_g197 (.A(G1464_285_gat), .Y(G5223_382_gat) );
AND2XL U_g198 (.A(G1501_291_gat), .B(G4442_290_gat), .Y(G2878_386_gat) );
AND2XL U_g199 (.A(G4514_292_gat), .B(G2857_293_gat), .Y(G2876_389_gat) );
AND2XL U_g200 (.A(G575_309_gat), .B(G1184_294_gat), .Y(G280_391_gat) );
INVXL U_g201 (.A(G446_393_gat), .Y(G1477_394_gat) );
BUFX20 U_g202 (.A(G1210_298_gat), .Y(G6554_396_gat) );
BUFX20 U_g203 (.A(G1210_298_gat), .Y(G6514_397_gat) );
BUFX20 U_g204 (.A(G1198_299_gat), .Y(G5186_398_gat) );
BUFX20 U_g205 (.A(G1198_299_gat), .Y(G5178_399_gat) );
BUFX20 U_g206 (.A(G1198_299_gat), .Y(G4916_400_gat) );
BUFX20 U_g207 (.A(G1198_299_gat), .Y(G4876_401_gat) );
BUFX20 U_g208 (.A(G1512_300_gat), .Y(G587_402_gat) );
BUFX20 U_g209 (.A(G1512_300_gat), .Y(G606_403_gat) );
BUFX20 U_g210 (.A(G1512_300_gat), .Y(G657_404_gat) );
BUFX20 U_g211 (.A(G1512_300_gat), .Y(G1336_405_gat) );
INVXL U_g212 (.A(G1512_300_gat), .Y(G1514_406_gat) );
BUFX20 U_g213 (.A(G1524_301_gat), .Y(G3622_407_gat) );
BUFX20 U_g214 (.A(G1524_301_gat), .Y(G3635_408_gat) );
BUFX20 U_g215 (.A(G1524_301_gat), .Y(G4640_409_gat) );
BUFX20 U_g216 (.A(G1524_301_gat), .Y(G4653_410_gat) );
INVXL U_g217 (.A(G1524_301_gat), .Y(G1530_411_gat) );
BUFX20 U_g218 (.A(G1535_302_gat), .Y(G3755_412_gat) );
BUFX20 U_g219 (.A(G1535_302_gat), .Y(G2259_413_gat) );
BUFX20 U_g220 (.A(G1503_303_gat), .Y(G678_414_gat) );
BUFX20 U_g221 (.A(G1503_303_gat), .Y(G1350_415_gat) );
BUFX20 U_g222 (.A(G1503_303_gat), .Y(G2892_416_gat) );
BUFX20 U_g223 (.A(G1503_303_gat), .Y(G2909_417_gat) );
INVXL U_g224 (.A(G1503_303_gat), .Y(G1507_418_gat) );
BUFX20 U_g225 (.A(G1206_306_gat), .Y(G581_421_gat) );
BUFX20 U_g226 (.A(G1206_306_gat), .Y(G601_422_gat) );
BUFX20 U_g227 (.A(G1206_306_gat), .Y(G650_423_gat) );
BUFX20 U_g228 (.A(G1207_307_gat), .Y(G671_424_gat) );
BUFX20 U_g229 (.A(G1207_307_gat), .Y(G2886_425_gat) );
BUFX20 U_g230 (.A(G1207_307_gat), .Y(G2905_426_gat) );
BUFX20 U_g231 (.A(G432_428_gat), .Y(G453_596_gat) );
BUFX20 U_g232 (.A(G2883_314_gat), .Y(G6511_429_gat) );
INVXL U_g233 (.A(G2871_315_gat), .Y(G2872_430_gat) );
INVXL U_g234 (.A(G6853_318_gat), .Y(G6859_431_gat) );
INVXL U_g235 (.A(G6567_319_gat), .Y(G6573_432_gat) );
INVXL U_g236 (.A(G6575_320_gat), .Y(G6581_433_gat) );
INVXL U_g237 (.A(G6861_321_gat), .Y(G6867_434_gat) );
INVXL U_g238 (.A(G6583_322_gat), .Y(G6589_435_gat) );
INVXL U_g239 (.A(G6869_323_gat), .Y(G6875_436_gat) );
INVXL U_g240 (.A(G6909_324_gat), .Y(G6915_437_gat) );
INVXL U_g241 (.A(G6591_325_gat), .Y(G6597_438_gat) );
INVXL U_g242 (.A(G6877_326_gat), .Y(G6883_439_gat) );
INVXL U_g243 (.A(G6599_327_gat), .Y(G6605_440_gat) );
INVXL U_g244 (.A(G6607_328_gat), .Y(G6613_441_gat) );
INVXL U_g245 (.A(G6885_329_gat), .Y(G6891_442_gat) );
INVXL U_g246 (.A(G6893_330_gat), .Y(G6899_443_gat) );
INVXL U_g247 (.A(G6615_331_gat), .Y(G6621_444_gat) );
INVXL U_g248 (.A(G6901_332_gat), .Y(G6907_445_gat) );
INVXL U_g249 (.A(G6623_333_gat), .Y(G6629_446_gat) );
INVXL U_g250 (.A(G6631_334_gat), .Y(G6637_447_gat) );
INVXL U_g251 (.A(G6917_335_gat), .Y(G6923_448_gat) );
INVXL U_g252 (.A(G5985_336_gat), .Y(G5991_449_gat) );
INVXL U_g253 (.A(G5865_337_gat), .Y(G5871_450_gat) );
INVXL U_g254 (.A(G5873_338_gat), .Y(G5879_451_gat) );
INVXL U_g255 (.A(G5993_339_gat), .Y(G5999_452_gat) );
INVXL U_g256 (.A(G6001_340_gat), .Y(G6007_453_gat) );
INVXL U_g257 (.A(G5881_341_gat), .Y(G5887_454_gat) );
INVXL U_g258 (.A(G6041_342_gat), .Y(G6047_455_gat) );
INVXL U_g259 (.A(G5889_343_gat), .Y(G5895_456_gat) );
INVXL U_g260 (.A(G5897_344_gat), .Y(G5903_457_gat) );
INVXL U_g261 (.A(G6009_345_gat), .Y(G6015_458_gat) );
INVXL U_g262 (.A(G6017_346_gat), .Y(G6023_459_gat) );
INVXL U_g263 (.A(G5905_347_gat), .Y(G5911_460_gat) );
INVXL U_g264 (.A(G5913_348_gat), .Y(G5919_461_gat) );
INVXL U_g265 (.A(G6025_349_gat), .Y(G6031_462_gat) );
INVXL U_g266 (.A(G6033_350_gat), .Y(G6039_463_gat) );
INVXL U_g267 (.A(G5921_351_gat), .Y(G5927_464_gat) );
AND2XL U_g268 (.A(G4653_410_gat), .B(G2258_249_gat), .Y(G4685_465_gat) );
INVXL U_g269 (.A(G5393_352_gat), .Y(G5399_466_gat) );
INVXL U_g270 (.A(G5745_353_gat), .Y(G5751_467_gat) );
AND2XL U_g271 (.A(G4653_410_gat), .B(G2255_252_gat), .Y(G4683_468_gat) );
INVXL U_g272 (.A(G5753_354_gat), .Y(G5759_469_gat) );
INVXL U_g273 (.A(G5401_355_gat), .Y(G5407_470_gat) );
AND2XL U_g274 (.A(G4653_410_gat), .B(G2249_255_gat), .Y(G4681_471_gat) );
INVXL U_g275 (.A(G5409_356_gat), .Y(G5415_472_gat) );
INVXL U_g276 (.A(G5761_357_gat), .Y(G5767_473_gat) );
INVXL U_g277 (.A(G5769_358_gat), .Y(G5775_474_gat) );
INVXL U_g278 (.A(G5449_359_gat), .Y(G5455_475_gat) );
AND2XL U_g279 (.A(G4653_410_gat), .B(G2241_257_gat), .Y(G4679_476_gat) );
AND2XL U_g280 (.A(G4653_410_gat), .B(G2238_259_gat), .Y(G4677_477_gat) );
INVXL U_g281 (.A(G5417_360_gat), .Y(G5423_478_gat) );
INVXL U_g282 (.A(G5777_361_gat), .Y(G5783_479_gat) );
INVXL U_g283 (.A(G5785_362_gat), .Y(G5791_480_gat) );
INVXL U_g284 (.A(G5425_363_gat), .Y(G5431_481_gat) );
AND2XL U_g285 (.A(G4640_409_gat), .B(G2232_262_gat), .Y(G4675_482_gat) );
AND2XL U_g286 (.A(G4640_409_gat), .B(G2226_264_gat), .Y(G4673_483_gat) );
INVXL U_g287 (.A(G5433_364_gat), .Y(G5439_484_gat) );
INVXL U_g288 (.A(G5793_365_gat), .Y(G5799_485_gat) );
INVXL U_g289 (.A(G5801_366_gat), .Y(G5807_486_gat) );
INVXL U_g290 (.A(G5441_367_gat), .Y(G5447_487_gat) );
AND2XL U_g291 (.A(G4640_409_gat), .B(G2220_266_gat), .Y(G4671_488_gat) );
INVXL U_g292 (.A(G5457_368_gat), .Y(G5463_489_gat) );
AND2XL U_g293 (.A(G4640_409_gat), .B(G2213_268_gat), .Y(G4669_490_gat) );
INVXL U_g294 (.A(G5809_369_gat), .Y(G5815_491_gat) );
AND2XL U_g295 (.A(G4640_409_gat), .B(G2210_270_gat), .Y(G4667_492_gat) );
AND2XL U_g296 (.A(G3635_408_gat), .B(G1499_273_gat), .Y(G3663_493_gat) );
INVXL U_g297 (.A(G5175_372_gat), .Y(G5181_494_gat) );
INVXL U_g298 (.A(G4873_373_gat), .Y(G4879_495_gat) );
AND2XL U_g299 (.A(G3635_408_gat), .B(G1495_276_gat), .Y(G3661_496_gat) );
BUFX20 U_g300 (.A(G1519_374_gat), .Y(G4913_497_gat) );
BUFX20 U_g301 (.A(G1519_374_gat), .Y(G5183_498_gat) );
AND2XL U_g302 (.A(G3635_408_gat), .B(G1488_279_gat), .Y(G3659_499_gat) );
INVXL U_g303 (.A(G4881_375_gat), .Y(G4887_500_gat) );
INVXL U_g304 (.A(G5191_376_gat), .Y(G5197_501_gat) );
INVXL U_g305 (.A(G5199_377_gat), .Y(G5205_502_gat) );
INVXL U_g306 (.A(G4889_378_gat), .Y(G4895_503_gat) );
AND2XL U_g307 (.A(G3622_407_gat), .B(G1482_281_gat), .Y(G3657_504_gat) );
INVXL U_g308 (.A(G5215_379_gat), .Y(G5221_505_gat) );
AND2XL U_g309 (.A(G3622_407_gat), .B(G1471_283_gat), .Y(G3653_506_gat) );
INVXL U_g310 (.A(G4905_380_gat), .Y(G4911_507_gat) );
INVXL U_g311 (.A(G4921_381_gat), .Y(G4927_508_gat) );
AND2XL U_g312 (.A(G3622_407_gat), .B(G1464_285_gat), .Y(G3651_509_gat) );
INVXL U_g313 (.A(G5223_382_gat), .Y(G5229_510_gat) );
AND2XL U_g314 (.A(G3622_407_gat), .B(G1461_287_gat), .Y(G3649_511_gat) );
AND2XL U_g315 (.A(G2892_416_gat), .B(G216_139_gat), .Y(G2921_512_gat) );
AND2XL U_g316 (.A(G2892_416_gat), .B(G215_138_gat), .Y(G2923_513_gat) );
AND2XL U_g317 (.A(G2892_416_gat), .B(G214_137_gat), .Y(G2925_514_gat) );
AND2XL U_g318 (.A(G2909_417_gat), .B(G213_136_gat), .Y(G2927_515_gat) );
AND2XL U_g319 (.A(G2909_417_gat), .B(G212_135_gat), .Y(G2929_516_gat) );
AND2XL U_g320 (.A(G2909_417_gat), .B(G211_134_gat), .Y(G2931_517_gat) );
AND2XL U_g321 (.A(G2892_416_gat), .B(G209_132_gat), .Y(G2919_518_gat) );
AND2XL U_g322 (.A(G1336_405_gat), .B(G181_104_gat), .Y(G1364_519_gat) );
AND2XL U_g323 (.A(G1336_405_gat), .B(G180_103_gat), .Y(G1368_520_gat) );
AND2XL U_g324 (.A(G1336_405_gat), .B(G179_102_gat), .Y(G1370_521_gat) );
AND2XL U_g325 (.A(G1336_405_gat), .B(G178_101_gat), .Y(G1372_522_gat) );
AND2XL U_g326 (.A(G657_404_gat), .B(G177_100_gat), .Y(G691_523_gat) );
AND2XL U_g327 (.A(G657_404_gat), .B(G176_99_gat), .Y(G693_524_gat) );
AND2XL U_g328 (.A(G657_404_gat), .B(G175_98_gat), .Y(G695_525_gat) );
AND2XL U_g329 (.A(G657_404_gat), .B(G174_97_gat), .Y(G697_526_gat) );
AND2XL U_g330 (.A(G657_404_gat), .B(G173_96_gat), .Y(G699_527_gat) );
AND2XL U_g331 (.A(G1336_405_gat), .B(G171_94_gat), .Y(G1366_528_gat) );
AND2XL U_g332 (.A(G587_402_gat), .B(G170_93_gat), .Y(G615_529_gat) );
AND2XL U_g333 (.A(G587_402_gat), .B(G169_92_gat), .Y(G617_530_gat) );
AND2XL U_g334 (.A(G587_402_gat), .B(G168_91_gat), .Y(G619_531_gat) );
AND2XL U_g335 (.A(G587_402_gat), .B(G167_90_gat), .Y(G621_532_gat) );
AND2XL U_g336 (.A(G606_403_gat), .B(G166_89_gat), .Y(G623_533_gat) );
AND2XL U_g337 (.A(G606_403_gat), .B(G165_88_gat), .Y(G625_534_gat) );
AND2XL U_g338 (.A(G606_403_gat), .B(G164_87_gat), .Y(G627_535_gat) );
AND2XL U_g339 (.A(G1350_415_gat), .B(G161_84_gat), .Y(G1374_537_gat) );
AND2XL U_g340 (.A(G1350_415_gat), .B(G160_83_gat), .Y(G1378_538_gat) );
AND2XL U_g341 (.A(G1350_415_gat), .B(G159_82_gat), .Y(G1380_539_gat) );
AND2XL U_g342 (.A(G1350_415_gat), .B(G158_81_gat), .Y(G1382_540_gat) );
AND2XL U_g343 (.A(G678_414_gat), .B(G157_80_gat), .Y(G701_541_gat) );
AND2XL U_g344 (.A(G678_414_gat), .B(G156_79_gat), .Y(G703_542_gat) );
AND2XL U_g345 (.A(G678_414_gat), .B(G155_78_gat), .Y(G705_543_gat) );
AND2XL U_g346 (.A(G678_414_gat), .B(G154_77_gat), .Y(G707_544_gat) );
AND2XL U_g347 (.A(G678_414_gat), .B(G153_76_gat), .Y(G709_545_gat) );
AND2XL U_g348 (.A(G1350_415_gat), .B(G151_74_gat), .Y(G1376_546_gat) );
BUFX20 U_g349 (.A(G1477_394_gat), .Y(G4897_548_gat) );
BUFX20 U_g350 (.A(G1477_394_gat), .Y(G5207_549_gat) );
AND2XL U_g351 (.A(G3622_407_gat), .B(G1500_296_gat), .Y(G3655_550_gat) );
AND2XL U_g352 (.A(G3755_412_gat), .B(G66_29_gat), .Y(G3790_551_gat) );
AND2XL U_g353 (.A(G3755_412_gat), .B(G50_15_gat), .Y(G3788_552_gat) );
AND2XL U_g354 (.A(G3755_412_gat), .B(G47_14_gat), .Y(G3782_553_gat) );
AND2XL U_g355 (.A(G2259_413_gat), .B(G44_13_gat), .Y(G2286_554_gat) );
AND2XL U_g356 (.A(G2259_413_gat), .B(G41_12_gat), .Y(G2288_555_gat) );
INVXL U_g357 (.A(G6554_396_gat), .Y(G6558_556_gat) );
AND2XL U_g358 (.A(G1210_298_gat), .B(G2883_314_gat), .Y(G3221_557_gat) );
INVXL U_g359 (.A(G6514_397_gat), .Y(G6518_558_gat) );
AND2XL U_g360 (.A(G1198_299_gat), .B(G1519_374_gat), .Y(G784_559_gat) );
AND2XL U_g361 (.A(G1519_374_gat), .B(G1198_299_gat), .Y(G1014_560_gat) );
AND2XL U_g362 (.A(G1519_374_ngat), .B(G1198_299_ngat), .Y(G5231_561_gat) );
INVXL U_g363 (.A(G5186_398_gat), .Y(G5190_562_gat) );
INVXL U_g364 (.A(G5178_399_gat), .Y(G5182_563_gat) );
AND2XL U_g365 (.A(G1198_299_ngat), .B(G1519_374_ngat), .Y(G4929_564_gat) );
INVXL U_g366 (.A(G4916_400_gat), .Y(G4920_565_gat) );
INVXL U_g367 (.A(G4876_401_gat), .Y(G4880_566_gat) );
AND2XL U_g368 (.A(G3755_412_gat), .B(G35_10_gat), .Y(G3784_567_gat) );
AND2XL U_g369 (.A(G3755_412_gat), .B(G32_9_gat), .Y(G3786_568_gat) );
AND2XL U_g370 (.A(G2259_413_gat), .B(G29_8_gat), .Y(G2290_569_gat) );
AND2XL U_g371 (.A(G2259_413_gat), .B(G26_7_gat), .Y(G2292_570_gat) );
AND2XL U_g372 (.A(G2259_413_gat), .B(G23_6_gat), .Y(G2294_571_gat) );
INVXL U_g373 (.A(G587_402_gat), .Y(G594_572_gat) );
INVXL U_g374 (.A(G606_403_gat), .Y(G611_573_gat) );
INVXL U_g375 (.A(G657_404_gat), .Y(G664_574_gat) );
INVXL U_g376 (.A(G1336_405_gat), .Y(G1343_575_gat) );
BUFX20 U_g377 (.A(G1514_406_gat), .Y(G2019_576_gat) );
BUFX20 U_g378 (.A(G1514_406_gat), .Y(G2117_577_gat) );
INVXL U_g379 (.A(G3622_407_gat), .Y(G3629_578_gat) );
INVXL U_g380 (.A(G3635_408_gat), .Y(G3642_579_gat) );
INVXL U_g381 (.A(G4640_409_gat), .Y(G4647_580_gat) );
INVXL U_g382 (.A(G4653_410_gat), .Y(G4660_581_gat) );
BUFX20 U_g383 (.A(G1530_411_gat), .Y(G4444_582_gat) );
BUFX20 U_g384 (.A(G1530_411_gat), .Y(G4457_583_gat) );
BUFX20 U_g385 (.A(G1530_411_gat), .Y(G4094_584_gat) );
BUFX20 U_g386 (.A(G1530_411_gat), .Y(G4107_585_gat) );
INVXL U_g387 (.A(G3755_412_gat), .Y(G3762_586_gat) );
INVXL U_g388 (.A(G2259_413_gat), .Y(G2266_587_gat) );
INVXL U_g389 (.A(G678_414_gat), .Y(G685_588_gat) );
INVXL U_g390 (.A(G1350_415_gat), .Y(G1357_589_gat) );
INVXL U_g391 (.A(G2892_416_gat), .Y(G2899_590_gat) );
INVXL U_g392 (.A(G2909_417_gat), .Y(G2914_591_gat) );
BUFX20 U_g393 (.A(G1507_418_gat), .Y(G2032_592_gat) );
BUFX20 U_g394 (.A(G1507_418_gat), .Y(G2130_593_gat) );
BUFX20 U_g395 (.A(G1507_418_gat), .Y(G2272_594_gat) );
BUFX20 U_g396 (.A(G1507_418_gat), .Y(G3768_595_gat) );
OR2XL U_g397 (.A(G6518_558_ngat), .B(G6511_429_ngat), .Y(G3169_597_gat) );
INVXL U_g398 (.A(G6511_429_gat), .Y(G6517_598_gat) );
BUFX20 U_g399 (.A(G2872_430_gat), .Y(G6551_599_gat) );
AND2XL U_g400 (.A(G3642_579_gat), .B(G3703_245_gat), .Y(G3665_600_gat) );
AND2XL U_g401 (.A(G3642_579_gat), .B(G2204_174_gat), .Y(G3662_601_gat) );
OR2XL U_g402 (.A(G5182_563_ngat), .B(G5175_372_ngat), .Y(G1006_602_gat) );
OR2XL U_g403 (.A(G4880_566_ngat), .B(G4873_373_ngat), .Y(G764_603_gat) );
OR2XL U_g404 (.A(G4920_565_ngat), .B(G4913_497_ngat), .Y(G886_604_gat) );
INVXL U_g405 (.A(G4913_497_gat), .Y(G4919_605_gat) );
OR2XL U_g406 (.A(G5190_562_ngat), .B(G5183_498_ngat), .Y(G1018_606_gat) );
INVXL U_g407 (.A(G5183_498_gat), .Y(G5189_607_gat) );
AND2XL U_g408 (.A(G3642_579_gat), .B(G1455_166_gat), .Y(G3660_608_gat) );
OR2XL U_g409 (.A(G2921_512_gat), .B(G2899_590_gat), .Y(G2922_609_gat) );
OR2XL U_g410 (.A(G2923_513_gat), .B(G2899_590_gat), .Y(G2924_610_gat) );
OR2XL U_g411 (.A(G2925_514_gat), .B(G2899_590_gat), .Y(G2926_611_gat) );
OR2XL U_g412 (.A(G2927_515_gat), .B(G2914_591_gat), .Y(G2928_612_gat) );
OR2XL U_g413 (.A(G2929_516_gat), .B(G2914_591_gat), .Y(G2930_613_gat) );
OR2XL U_g414 (.A(G2931_517_gat), .B(G2914_591_gat), .Y(G2932_614_gat) );
OR2XL U_g415 (.A(G2919_518_gat), .B(G2899_590_gat), .Y(G2920_615_gat) );
AND2XL U_g416 (.A(G2266_587_gat), .B(G208_131_gat), .Y(G2285_616_gat) );
AND2XL U_g417 (.A(G2266_587_gat), .B(G207_130_gat), .Y(G2289_617_gat) );
AND2XL U_g418 (.A(G2266_587_gat), .B(G206_129_gat), .Y(G2291_618_gat) );
AND2XL U_g419 (.A(G2266_587_gat), .B(G205_128_gat), .Y(G2293_619_gat) );
AND2XL U_g420 (.A(G2266_587_gat), .B(G198_121_gat), .Y(G2287_620_gat) );
AND2XL U_g421 (.A(G3762_586_gat), .B(G193_116_gat), .Y(G3781_621_gat) );
AND2XL U_g422 (.A(G3762_586_gat), .B(G192_115_gat), .Y(G3783_622_gat) );
AND2XL U_g423 (.A(G3762_586_gat), .B(G191_114_gat), .Y(G3785_623_gat) );
AND2XL U_g424 (.A(G3762_586_gat), .B(G190_113_gat), .Y(G3787_624_gat) );
AND2XL U_g425 (.A(G3762_586_gat), .B(G189_112_gat), .Y(G3789_625_gat) );
OR2XL U_g426 (.A(G691_523_gat), .B(G664_574_gat), .Y(G692_626_gat) );
OR2XL U_g427 (.A(G693_524_gat), .B(G664_574_gat), .Y(G694_627_gat) );
OR2XL U_g428 (.A(G695_525_gat), .B(G664_574_gat), .Y(G696_628_gat) );
OR2XL U_g429 (.A(G697_526_gat), .B(G664_574_gat), .Y(G698_629_gat) );
OR2XL U_g430 (.A(G699_527_gat), .B(G664_574_gat), .Y(G700_630_gat) );
OR2XL U_g431 (.A(G615_529_gat), .B(G594_572_gat), .Y(G577_631_gat) );
OR2XL U_g432 (.A(G617_530_gat), .B(G594_572_gat), .Y(G618_632_gat) );
OR2XL U_g433 (.A(G619_531_gat), .B(G594_572_gat), .Y(G620_633_gat) );
OR2XL U_g434 (.A(G621_532_gat), .B(G594_572_gat), .Y(G622_634_gat) );
OR2XL U_g435 (.A(G623_533_gat), .B(G611_573_gat), .Y(G624_635_gat) );
OR2XL U_g436 (.A(G625_534_gat), .B(G611_573_gat), .Y(G626_636_gat) );
OR2XL U_g437 (.A(G627_535_gat), .B(G611_573_gat), .Y(G628_637_gat) );
OR2XL U_g438 (.A(G701_541_gat), .B(G685_588_gat), .Y(G702_638_gat) );
OR2XL U_g439 (.A(G703_542_gat), .B(G685_588_gat), .Y(G704_639_gat) );
OR2XL U_g440 (.A(G705_543_gat), .B(G685_588_gat), .Y(G706_640_gat) );
OR2XL U_g441 (.A(G707_544_gat), .B(G685_588_gat), .Y(G708_641_gat) );
OR2XL U_g442 (.A(G709_545_gat), .B(G685_588_gat), .Y(G710_642_gat) );
AND2XL U_g443 (.A(G1357_589_gat), .B(G147_72_gat), .Y(G1375_643_gat) );
AND2XL U_g444 (.A(G1343_575_gat), .B(G147_72_gat), .Y(G1365_644_gat) );
AND2XL U_g445 (.A(G1357_589_gat), .B(G144_71_gat), .Y(G1379_645_gat) );
AND2XL U_g446 (.A(G1343_575_gat), .B(G144_71_gat), .Y(G1369_646_gat) );
AND2XL U_g447 (.A(G1343_575_gat), .B(G141_70_gat), .Y(G1363_647_gat) );
AND2XL U_g448 (.A(G1357_589_gat), .B(G141_70_gat), .Y(G1373_648_gat) );
AND2XL U_g449 (.A(G1357_589_gat), .B(G138_69_gat), .Y(G1377_649_gat) );
AND2XL U_g450 (.A(G1343_575_gat), .B(G138_69_gat), .Y(G1367_650_gat) );
AND2XL U_g451 (.A(G1357_589_gat), .B(G135_68_gat), .Y(G1381_651_gat) );
AND2XL U_g452 (.A(G1343_575_gat), .B(G135_68_gat), .Y(G1371_652_gat) );
AND2XL U_g453 (.A(G2019_576_gat), .B(G130_65_gat), .Y(G2048_653_gat) );
AND2XL U_g454 (.A(G2032_592_gat), .B(G130_65_gat), .Y(G2058_654_gat) );
AND2XL U_g455 (.A(G2032_592_gat), .B(G127_64_gat), .Y(G2060_655_gat) );
AND2XL U_g456 (.A(G2019_576_gat), .B(G127_64_gat), .Y(G2050_656_gat) );
AND2XL U_g457 (.A(G2032_592_gat), .B(G124_63_gat), .Y(G2062_657_gat) );
AND2XL U_g458 (.A(G2019_576_gat), .B(G124_63_gat), .Y(G2052_658_gat) );
AND2XL U_g459 (.A(G2130_593_gat), .B(G121_62_gat), .Y(G2162_659_gat) );
AND2XL U_g460 (.A(G2117_577_gat), .B(G121_62_gat), .Y(G2152_660_gat) );
AND2XL U_g461 (.A(G2117_577_gat), .B(G118_61_gat), .Y(G2146_661_gat) );
AND2XL U_g462 (.A(G2130_593_gat), .B(G118_61_gat), .Y(G2156_662_gat) );
AND2XL U_g463 (.A(G2117_577_gat), .B(G115_60_gat), .Y(G2144_663_gat) );
AND2XL U_g464 (.A(G2130_593_gat), .B(G115_60_gat), .Y(G2154_664_gat) );
AND2XL U_g465 (.A(G3629_578_gat), .B(G114_59_gat), .Y(G3648_665_gat) );
AND2XL U_g466 (.A(G3629_578_gat), .B(G113_58_gat), .Y(G3650_666_gat) );
AND2XL U_g467 (.A(G3629_578_gat), .B(G112_57_gat), .Y(G3656_667_gat) );
AND2XL U_g468 (.A(G3629_578_gat), .B(G111_56_gat), .Y(G3652_668_gat) );
AND2XL U_g469 (.A(G4660_581_gat), .B(G110_55_gat), .Y(G4684_669_gat) );
AND2XL U_g470 (.A(G4660_581_gat), .B(G109_54_gat), .Y(G4682_670_gat) );
INVXL U_g471 (.A(G4897_548_gat), .Y(G4903_671_gat) );
INVXL U_g472 (.A(G5207_549_gat), .Y(G5213_672_gat) );
AND2XL U_g473 (.A(G2019_576_gat), .B(G103_52_gat), .Y(G2046_673_gat) );
AND2XL U_g474 (.A(G2032_592_gat), .B(G103_52_gat), .Y(G2056_674_gat) );
AND2XL U_g475 (.A(G2032_592_gat), .B(G100_51_gat), .Y(G2064_675_gat) );
AND2XL U_g476 (.A(G2019_576_gat), .B(G100_51_gat), .Y(G2054_676_gat) );
AND2XL U_g477 (.A(G2130_593_gat), .B(G97_50_gat), .Y(G2158_677_gat) );
AND2XL U_g478 (.A(G2117_577_gat), .B(G97_50_gat), .Y(G2148_678_gat) );
AND2XL U_g479 (.A(G2130_593_gat), .B(G94_49_gat), .Y(G2160_679_gat) );
AND2XL U_g480 (.A(G2117_577_gat), .B(G94_49_gat), .Y(G2150_680_gat) );
AND2XL U_g481 (.A(G3642_579_gat), .B(G88_47_gat), .Y(G3658_681_gat) );
AND2XL U_g482 (.A(G3629_578_gat), .B(G87_46_gat), .Y(G3654_682_gat) );
AND2XL U_g483 (.A(G4660_581_gat), .B(G86_45_gat), .Y(G4680_683_gat) );
AND2XL U_g484 (.A(G4647_580_gat), .B(G85_44_gat), .Y(G4674_684_gat) );
AND2XL U_g485 (.A(G4647_580_gat), .B(G84_43_gat), .Y(G4672_685_gat) );
AND2XL U_g486 (.A(G4647_580_gat), .B(G83_42_gat), .Y(G4670_686_gat) );
AND2XL U_g487 (.A(G4647_580_gat), .B(G82_41_gat), .Y(G4666_687_gat) );
AND2XL U_g488 (.A(G4094_584_gat), .B(G81_40_gat), .Y(G4135_688_gat) );
AND2XL U_g489 (.A(G4107_585_gat), .B(G80_39_gat), .Y(G4138_689_gat) );
AND2XL U_g490 (.A(G4107_585_gat), .B(G79_38_gat), .Y(G4141_690_gat) );
AND2XL U_g491 (.A(G4094_584_gat), .B(G78_37_gat), .Y(G4129_691_gat) );
AND2XL U_g492 (.A(G4094_584_gat), .B(G77_36_gat), .Y(G4126_692_gat) );
AND2XL U_g493 (.A(G4444_582_gat), .B(G76_35_gat), .Y(G4477_693_gat) );
AND2XL U_g494 (.A(G4444_582_gat), .B(G75_34_gat), .Y(G4479_694_gat) );
AND2XL U_g495 (.A(G4444_582_gat), .B(G74_33_gat), .Y(G4475_695_gat) );
AND2XL U_g496 (.A(G4457_583_gat), .B(G73_32_gat), .Y(G4481_696_gat) );
AND2XL U_g497 (.A(G4444_582_gat), .B(G70_31_gat), .Y(G4473_697_gat) );
AND2XL U_g498 (.A(G3642_579_gat), .B(G70_31_gat), .Y(G3666_698_gat) );
AND2XL U_g499 (.A(G4444_582_gat), .B(G69_30_gat), .Y(G4471_699_gat) );
AND2XL U_g500 (.A(G3768_595_gat), .B(G66_29_gat), .Y(G3800_700_gat) );
AND2XL U_g501 (.A(G4647_580_gat), .B(G65_28_gat), .Y(G4668_701_gat) );
AND2XL U_g502 (.A(G4660_581_gat), .B(G64_27_gat), .Y(G4676_702_gat) );
AND2XL U_g503 (.A(G4660_581_gat), .B(G63_26_gat), .Y(G4678_703_gat) );
AND2XL U_g504 (.A(G4107_585_gat), .B(G62_25_gat), .Y(G4150_704_gat) );
AND2XL U_g505 (.A(G4107_585_gat), .B(G61_24_gat), .Y(G4147_705_gat) );
AND2XL U_g506 (.A(G4107_585_gat), .B(G60_23_gat), .Y(G4144_706_gat) );
AND2XL U_g507 (.A(G4094_584_gat), .B(G59_22_gat), .Y(G4132_707_gat) );
AND2XL U_g508 (.A(G4094_584_gat), .B(G58_21_gat), .Y(G4123_708_gat) );
AND2XL U_g509 (.A(G4457_583_gat), .B(G56_19_gat), .Y(G4489_709_gat) );
AND2XL U_g510 (.A(G4457_583_gat), .B(G55_18_gat), .Y(G4487_710_gat) );
AND2XL U_g511 (.A(G4457_583_gat), .B(G54_17_gat), .Y(G4485_711_gat) );
AND2XL U_g512 (.A(G4457_583_gat), .B(G53_16_gat), .Y(G4483_712_gat) );
AND2XL U_g513 (.A(G3768_595_gat), .B(G50_15_gat), .Y(G3798_713_gat) );
AND2XL U_g514 (.A(G3768_595_gat), .B(G47_14_gat), .Y(G3792_714_gat) );
AND2XL U_g515 (.A(G2272_594_gat), .B(G44_13_gat), .Y(G2296_715_gat) );
AND2XL U_g516 (.A(G2272_594_gat), .B(G41_12_gat), .Y(G2298_716_gat) );
AND2XL U_g517 (.A(G1210_298_gat), .B(G2872_430_gat), .Y(G3173_717_gat) );
BUFX20 U_g518 (.A(G784_559_gat), .Y(G4970_718_gat) );
BUFX20 U_g519 (.A(G1014_560_gat), .Y(G5239_719_gat) );
INVXL U_g520 (.A(G5231_561_gat), .Y(G5237_720_gat) );
OR2XL U_g521 (.A(G5181_494_ngat), .B(G5178_399_ngat), .Y(G1005_721_gat) );
INVXL U_g522 (.A(G4929_564_gat), .Y(G4935_722_gat) );
OR2XL U_g523 (.A(G4879_495_ngat), .B(G4876_401_ngat), .Y(G763_723_gat) );
AND2XL U_g524 (.A(G3768_595_gat), .B(G35_10_gat), .Y(G3794_724_gat) );
AND2XL U_g525 (.A(G3768_595_gat), .B(G32_9_gat), .Y(G3796_725_gat) );
AND2XL U_g526 (.A(G2272_594_gat), .B(G29_8_gat), .Y(G2300_726_gat) );
AND2XL U_g527 (.A(G2272_594_gat), .B(G26_7_gat), .Y(G2302_727_gat) );
AND2XL U_g528 (.A(G2272_594_gat), .B(G23_6_gat), .Y(G2304_728_gat) );
OR2XL U_g529 (.A(G587_402_gat), .B(G594_572_gat), .Y(G616_729_gat) );
INVXL U_g530 (.A(G2019_576_gat), .Y(G2026_730_gat) );
INVXL U_g531 (.A(G2117_577_gat), .Y(G2124_731_gat) );
INVXL U_g532 (.A(G4444_582_gat), .Y(G4451_732_gat) );
INVXL U_g533 (.A(G4457_583_gat), .Y(G4464_733_gat) );
INVXL U_g534 (.A(G4094_584_gat), .Y(G4101_734_gat) );
INVXL U_g535 (.A(G4107_585_gat), .Y(G4114_735_gat) );
OR2XL U_g536 (.A(G2892_416_gat), .B(G2899_590_gat), .Y(G2918_736_gat) );
INVXL U_g537 (.A(G2032_592_gat), .Y(G2039_737_gat) );
INVXL U_g538 (.A(G2130_593_gat), .Y(G2137_738_gat) );
INVXL U_g539 (.A(G2272_594_gat), .Y(G2279_739_gat) );
INVXL U_g540 (.A(G3768_595_gat), .Y(G3775_740_gat) );
INVXL U_g541 (.A(G6551_599_gat), .Y(G6557_741_gat) );
AND2XL U_g542 (.A(G4114_735_gat), .B(G4439_209_gat), .Y(G4149_742_gat) );
AND2XL U_g543 (.A(G4114_735_gat), .B(G4434_211_gat), .Y(G4146_743_gat) );
AND2XL U_g544 (.A(G4114_735_gat), .B(G4429_213_gat), .Y(G4143_744_gat) );
AND2XL U_g545 (.A(G4114_735_gat), .B(G4422_215_gat), .Y(G4140_745_gat) );
AND2XL U_g546 (.A(G4114_735_gat), .B(G4417_217_gat), .Y(G4137_746_gat) );
AND2XL U_g547 (.A(G4101_734_gat), .B(G4412_219_gat), .Y(G4134_747_gat) );
AND2XL U_g548 (.A(G4101_734_gat), .B(G4407_221_gat), .Y(G4131_748_gat) );
AND2XL U_g549 (.A(G4101_734_gat), .B(G4402_223_gat), .Y(G4128_749_gat) );
AND2XL U_g550 (.A(G4101_734_gat), .B(G4396_225_gat), .Y(G4125_750_gat) );
AND2XL U_g551 (.A(G4101_734_gat), .B(G4121_228_gat), .Y(G4122_751_gat) );
AND2XL U_g552 (.A(G4464_733_gat), .B(G3751_229_gat), .Y(G4488_752_gat) );
AND2XL U_g553 (.A(G4464_733_gat), .B(G3745_231_gat), .Y(G4486_753_gat) );
AND2XL U_g554 (.A(G4464_733_gat), .B(G3739_233_gat), .Y(G4484_754_gat) );
AND2XL U_g555 (.A(G4464_733_gat), .B(G3731_235_gat), .Y(G4482_755_gat) );
AND2XL U_g556 (.A(G4464_733_gat), .B(G3725_237_gat), .Y(G4480_756_gat) );
AND2XL U_g557 (.A(G4451_732_gat), .B(G3719_239_gat), .Y(G4478_757_gat) );
AND2XL U_g558 (.A(G4451_732_gat), .B(G3713_241_gat), .Y(G4476_758_gat) );
AND2XL U_g559 (.A(G4451_732_gat), .B(G3707_243_gat), .Y(G4474_759_gat) );
AND2XL U_g560 (.A(G4451_732_gat), .B(G3703_245_gat), .Y(G4472_760_gat) );
AND2XL U_g561 (.A(G4451_732_gat), .B(G3700_247_gat), .Y(G4470_761_gat) );
OR2XL U_g562 (.A(G4685_465_gat), .B(G4684_669_gat), .Y(G4710_762_gat) );
OR2XL U_g563 (.A(G4683_468_gat), .B(G4682_670_gat), .Y(G4707_763_gat) );
OR2XL U_g564 (.A(G4681_471_gat), .B(G4680_683_gat), .Y(G4704_764_gat) );
OR2XL U_g565 (.A(G4679_476_gat), .B(G4678_703_gat), .Y(G4701_765_gat) );
OR2XL U_g566 (.A(G4677_477_gat), .B(G4676_702_gat), .Y(G4698_766_gat) );
OR2XL U_g567 (.A(G4675_482_gat), .B(G4674_684_gat), .Y(G4695_767_gat) );
OR2XL U_g568 (.A(G4673_483_gat), .B(G4672_685_gat), .Y(G4692_768_gat) );
OR2XL U_g569 (.A(G4671_488_gat), .B(G4670_686_gat), .Y(G4689_769_gat) );
OR2XL U_g570 (.A(G4669_490_gat), .B(G4668_701_gat), .Y(G4686_770_gat) );
OR2XL U_g571 (.A(G4667_492_gat), .B(G4666_687_gat), .Y(G7466_771_gat) );
OR2XL U_g572 (.A(G3663_493_gat), .B(G3662_601_gat), .Y(G6711_772_gat) );
OR2XL U_g573 (.A(G1006_602_ngat), .B(G1005_721_ngat), .Y(G1007_773_gat) );
OR2XL U_g574 (.A(G764_603_ngat), .B(G763_723_ngat), .Y(G765_774_gat) );
OR2XL U_g575 (.A(G3661_496_gat), .B(G3660_608_gat), .Y(G6714_775_gat) );
OR2XL U_g576 (.A(G3659_499_gat), .B(G3658_681_gat), .Y(G3679_776_gat) );
OR2XL U_g577 (.A(G3657_504_gat), .B(G3656_667_gat), .Y(G3676_777_gat) );
OR2XL U_g578 (.A(G3653_506_gat), .B(G3652_668_gat), .Y(G3670_778_gat) );
OR2XL U_g579 (.A(G3651_509_gat), .B(G3650_666_gat), .Y(G3667_779_gat) );
OR2XL U_g580 (.A(G3649_511_gat), .B(G3648_665_gat), .Y(G6690_780_gat) );
AND2XL U_g581 (.A(G2279_739_gat), .B(G239_162_gat), .Y(G2295_781_gat) );
AND2XL U_g582 (.A(G2279_739_gat), .B(G238_161_gat), .Y(G2299_782_gat) );
AND2XL U_g583 (.A(G2279_739_gat), .B(G237_160_gat), .Y(G2301_783_gat) );
AND2XL U_g584 (.A(G2279_739_gat), .B(G236_159_gat), .Y(G2303_784_gat) );
AND2XL U_g585 (.A(G2039_737_gat), .B(G235_158_gat), .Y(G2055_785_gat) );
AND2XL U_g586 (.A(G2039_737_gat), .B(G234_157_gat), .Y(G2057_786_gat) );
AND2XL U_g587 (.A(G2039_737_gat), .B(G233_156_gat), .Y(G2059_787_gat) );
AND2XL U_g588 (.A(G2039_737_gat), .B(G232_155_gat), .Y(G2061_788_gat) );
AND2XL U_g589 (.A(G2039_737_gat), .B(G231_154_gat), .Y(G2063_789_gat) );
AND2XL U_g590 (.A(G2279_739_gat), .B(G229_152_gat), .Y(G2297_790_gat) );
AND2XL U_g591 (.A(G2137_738_gat), .B(G227_150_gat), .Y(G2153_791_gat) );
AND2XL U_g592 (.A(G2137_738_gat), .B(G226_149_gat), .Y(G2157_792_gat) );
AND2XL U_g593 (.A(G2137_738_gat), .B(G225_148_gat), .Y(G2159_793_gat) );
AND2XL U_g594 (.A(G2137_738_gat), .B(G224_147_gat), .Y(G2161_794_gat) );
AND2XL U_g595 (.A(G3775_740_gat), .B(G223_146_gat), .Y(G3791_795_gat) );
AND2XL U_g596 (.A(G3775_740_gat), .B(G222_145_gat), .Y(G3793_796_gat) );
AND2XL U_g597 (.A(G3775_740_gat), .B(G221_144_gat), .Y(G3795_797_gat) );
AND2XL U_g598 (.A(G3775_740_gat), .B(G220_143_gat), .Y(G3797_798_gat) );
AND2XL U_g599 (.A(G3775_740_gat), .B(G219_142_gat), .Y(G3799_799_gat) );
AND2XL U_g600 (.A(G2137_738_gat), .B(G217_140_gat), .Y(G2155_800_gat) );
AND2XL U_g601 (.A(G2026_730_gat), .B(G204_127_gat), .Y(G2045_801_gat) );
AND2XL U_g602 (.A(G2026_730_gat), .B(G203_126_gat), .Y(G2047_802_gat) );
AND2XL U_g603 (.A(G2026_730_gat), .B(G202_125_gat), .Y(G2049_803_gat) );
AND2XL U_g604 (.A(G2026_730_gat), .B(G201_124_gat), .Y(G2051_804_gat) );
AND2XL U_g605 (.A(G2026_730_gat), .B(G200_123_gat), .Y(G2053_805_gat) );
AND2XL U_g606 (.A(G2124_731_gat), .B(G197_120_gat), .Y(G2143_806_gat) );
AND2XL U_g607 (.A(G2124_731_gat), .B(G196_119_gat), .Y(G2147_807_gat) );
AND2XL U_g608 (.A(G2124_731_gat), .B(G195_118_gat), .Y(G2149_808_gat) );
AND2XL U_g609 (.A(G2124_731_gat), .B(G194_117_gat), .Y(G2151_809_gat) );
AND2XL U_g610 (.A(G2124_731_gat), .B(G187_110_gat), .Y(G2145_810_gat) );
OR2XL U_g611 (.A(G1364_519_gat), .B(G1363_647_gat), .Y(G7296_811_gat) );
OR2XL U_g612 (.A(G1368_520_gat), .B(G1367_650_gat), .Y(G1387_812_gat) );
OR2XL U_g613 (.A(G1370_521_gat), .B(G1369_646_gat), .Y(G1391_813_gat) );
OR2XL U_g614 (.A(G1372_522_gat), .B(G1371_652_gat), .Y(G1395_814_gat) );
OR2XL U_g615 (.A(G1366_528_gat), .B(G1365_644_gat), .Y(G1383_815_gat) );
OR2XL U_g616 (.A(G1374_537_gat), .B(G1373_648_gat), .Y(G5318_816_gat) );
OR2XL U_g617 (.A(G1378_538_gat), .B(G1377_649_gat), .Y(G1406_817_gat) );
OR2XL U_g618 (.A(G1380_539_gat), .B(G1379_645_gat), .Y(G1412_818_gat) );
OR2XL U_g619 (.A(G1382_540_gat), .B(G1381_651_gat), .Y(G1418_819_gat) );
OR2XL U_g620 (.A(G1376_546_gat), .B(G1375_643_gat), .Y(G1399_820_gat) );
OR2XL U_g621 (.A(G3655_550_gat), .B(G3654_682_gat), .Y(G3673_821_gat) );
OR2XL U_g622 (.A(G3790_551_gat), .B(G3789_625_gat), .Y(G3813_822_gat) );
OR2XL U_g623 (.A(G3788_552_gat), .B(G3787_624_gat), .Y(G3810_823_gat) );
OR2XL U_g624 (.A(G3782_553_gat), .B(G3781_621_gat), .Y(G3801_824_gat) );
OR2XL U_g625 (.A(G2286_554_gat), .B(G2285_616_gat), .Y(G7252_825_gat) );
OR2XL U_g626 (.A(G2288_555_gat), .B(G2287_620_gat), .Y(G2305_826_gat) );
OR2XL U_g627 (.A(G6558_556_ngat), .B(G6551_599_ngat), .Y(G3211_827_gat) );
OR2XL U_g628 (.A(G6517_598_ngat), .B(G6514_397_ngat), .Y(G3168_828_gat) );
INVXL U_g629 (.A(G4970_718_gat), .Y(G4976_829_gat) );
INVXL U_g630 (.A(G5239_719_gat), .Y(G5245_830_gat) );
OR2XL U_g631 (.A(G5189_607_ngat), .B(G5186_398_ngat), .Y(G1017_831_gat) );
OR2XL U_g632 (.A(G4919_605_ngat), .B(G4916_400_ngat), .Y(G885_832_gat) );
OR2XL U_g633 (.A(G3784_567_gat), .B(G3783_622_gat), .Y(G3804_833_gat) );
OR2XL U_g634 (.A(G3786_568_gat), .B(G3785_623_gat), .Y(G3807_834_gat) );
OR2XL U_g635 (.A(G2290_569_gat), .B(G2289_617_gat), .Y(G2308_835_gat) );
OR2XL U_g636 (.A(G2292_570_gat), .B(G2291_618_gat), .Y(G2312_836_gat) );
OR2XL U_g637 (.A(G2294_571_gat), .B(G2293_619_gat), .Y(G2316_837_gat) );
OR2XL U_g638 (.A(G3635_408_gat), .B(G3666_698_gat), .Y(G3686_838_gat) );
OR2XL U_g639 (.A(G3635_408_gat), .B(G3665_600_gat), .Y(G3682_839_gat) );
AND2XL U_g640 (.A(G581_421_gat), .B(G577_631_gat), .Y(G579_840_gat) );
AND2XL U_g641 (.A(G581_421_gat), .B(G622_634_gat), .Y(G641_841_gat) );
AND2XL U_g642 (.A(G581_421_gat), .B(G620_633_gat), .Y(G637_842_gat) );
AND2XL U_g643 (.A(G581_421_gat), .B(G618_632_gat), .Y(G633_843_gat) );
AND2XL U_g644 (.A(G581_421_gat), .B(G616_729_gat), .Y(G629_844_gat) );
AND2XL U_g645 (.A(G601_422_gat), .B(G628_637_gat), .Y(G5305_845_gat) );
AND2XL U_g646 (.A(G601_422_gat), .B(G626_636_gat), .Y(G5308_846_gat) );
AND2XL U_g647 (.A(G601_422_gat), .B(G624_635_gat), .Y(G645_847_gat) );
AND2XL U_g648 (.A(G650_423_gat), .B(G700_630_gat), .Y(G727_848_gat) );
AND2XL U_g649 (.A(G650_423_gat), .B(G698_629_gat), .Y(G723_849_gat) );
AND2XL U_g650 (.A(G650_423_gat), .B(G696_628_gat), .Y(G719_850_gat) );
AND2XL U_g651 (.A(G650_423_gat), .B(G694_627_gat), .Y(G715_851_gat) );
AND2XL U_g652 (.A(G650_423_gat), .B(G692_626_gat), .Y(G711_852_gat) );
AND2XL U_g653 (.A(G671_424_gat), .B(G706_640_gat), .Y(G745_853_gat) );
AND2XL U_g654 (.A(G671_424_gat), .B(G704_639_gat), .Y(G737_854_gat) );
AND2XL U_g655 (.A(G671_424_gat), .B(G702_638_gat), .Y(G731_855_gat) );
AND2XL U_g656 (.A(G671_424_gat), .B(G710_642_gat), .Y(G757_856_gat) );
AND2XL U_g657 (.A(G671_424_gat), .B(G708_641_gat), .Y(G751_857_gat) );
AND2XL U_g658 (.A(G2886_425_gat), .B(G2926_611_gat), .Y(G2946_858_gat) );
AND2XL U_g659 (.A(G2886_425_gat), .B(G2924_610_gat), .Y(G2942_859_gat) );
AND2XL U_g660 (.A(G2886_425_gat), .B(G2922_609_gat), .Y(G2938_860_gat) );
AND2XL U_g661 (.A(G2886_425_gat), .B(G2920_615_gat), .Y(G2933_861_gat) );
AND2XL U_g662 (.A(G2886_425_gat), .B(G2918_736_gat), .Y(G4525_862_gat) );
AND2XL U_g663 (.A(G2905_426_gat), .B(G2932_614_gat), .Y(G5271_863_gat) );
AND2XL U_g664 (.A(G2905_426_gat), .B(G2930_613_gat), .Y(G5274_864_gat) );
AND2XL U_g665 (.A(G2905_426_gat), .B(G2928_612_gat), .Y(G2950_865_gat) );
OR2XL U_g666 (.A(G3169_597_ngat), .B(G3168_828_ngat), .Y(G3170_866_gat) );
AND2XL U_g667 (.A(G727_848_gat), .B(G4710_762_gat), .Y(G2962_867_gat) );
BUFX20 U_g668 (.A(G4710_762_gat), .Y(G7497_868_gat) );
BUFX20 U_g669 (.A(G4710_762_gat), .Y(G6367_869_gat) );
AND2XL U_g670 (.A(G757_856_gat), .B(G1192_251_gat), .Y(G1553_870_gat) );
AND2XL U_g671 (.A(G757_856_gat), .B(G1192_251_gat), .Y(G1802_871_gat) );
AND2XL U_g672 (.A(G723_849_gat), .B(G4707_763_gat), .Y(G2970_872_gat) );
BUFX20 U_g673 (.A(G4707_763_gat), .Y(G7500_873_gat) );
BUFX20 U_g674 (.A(G4707_763_gat), .Y(G6375_874_gat) );
AND2XL U_g675 (.A(G751_857_gat), .B(G1186_254_gat), .Y(G1816_875_gat) );
AND2XL U_g676 (.A(G751_857_gat), .B(G1186_254_gat), .Y(G1567_876_gat) );
AND2XL U_g677 (.A(G745_853_gat), .B(G2249_255_gat), .Y(G1584_877_gat) );
AND2XL U_g678 (.A(G745_853_gat), .B(G2249_255_gat), .Y(G1834_878_gat) );
AND2XL U_g679 (.A(G719_850_gat), .B(G4704_764_gat), .Y(G2977_879_gat) );
BUFX20 U_g680 (.A(G4704_764_gat), .Y(G6383_880_gat) );
BUFX20 U_g681 (.A(G4704_764_gat), .Y(G7487_881_gat) );
AND2XL U_g682 (.A(G737_854_gat), .B(G2241_257_gat), .Y(G1590_882_gat) );
AND2XL U_g683 (.A(G2241_257_gat), .B(G737_854_gat), .Y(G1841_883_gat) );
AND2XL U_g684 (.A(G2241_257_ngat), .B(G737_854_ngat), .Y(G5849_884_gat) );
AND2XL U_g685 (.A(G737_854_ngat), .B(G2241_257_ngat), .Y(G5465_885_gat) );
AND2XL U_g686 (.A(G715_851_gat), .B(G4701_765_gat), .Y(G2979_886_gat) );
BUFX20 U_g687 (.A(G4701_765_gat), .Y(G7490_887_gat) );
BUFX20 U_g688 (.A(G4701_765_gat), .Y(G6423_888_gat) );
AND2XL U_g689 (.A(G711_852_gat), .B(G4698_766_gat), .Y(G2989_889_gat) );
BUFX20 U_g690 (.A(G4698_766_gat), .Y(G7479_890_gat) );
BUFX20 U_g691 (.A(G4698_766_gat), .Y(G6391_891_gat) );
AND2XL U_g692 (.A(G731_855_gat), .B(G1178_261_gat), .Y(G1606_892_gat) );
AND2XL U_g693 (.A(G731_855_gat), .B(G1178_261_gat), .Y(G1866_893_gat) );
AND2XL U_g694 (.A(G1418_819_gat), .B(G2232_262_gat), .Y(G1624_894_gat) );
AND2XL U_g695 (.A(G1418_819_gat), .B(G2232_262_gat), .Y(G1880_895_gat) );
AND2XL U_g696 (.A(G1395_814_gat), .B(G4695_767_gat), .Y(G2998_896_gat) );
BUFX20 U_g697 (.A(G4695_767_gat), .Y(G6399_897_gat) );
BUFX20 U_g698 (.A(G4695_767_gat), .Y(G7482_898_gat) );
AND2XL U_g699 (.A(G1412_818_gat), .B(G2226_264_gat), .Y(G1647_899_gat) );
AND2XL U_g700 (.A(G1412_818_gat), .B(G2226_264_gat), .Y(G1897_900_gat) );
AND2XL U_g701 (.A(G1391_813_gat), .B(G4692_768_gat), .Y(G3006_901_gat) );
BUFX20 U_g702 (.A(G4692_768_gat), .Y(G7471_902_gat) );
BUFX20 U_g703 (.A(G4692_768_gat), .Y(G6407_903_gat) );
AND2XL U_g704 (.A(G1406_817_gat), .B(G2220_266_gat), .Y(G1669_904_gat) );
AND2XL U_g705 (.A(G1406_817_gat), .B(G2220_266_gat), .Y(G1914_905_gat) );
AND2XL U_g706 (.A(G1387_812_gat), .B(G4689_769_gat), .Y(G3013_906_gat) );
BUFX20 U_g707 (.A(G4689_769_gat), .Y(G6415_907_gat) );
BUFX20 U_g708 (.A(G4689_769_gat), .Y(G7474_908_gat) );
AND2XL U_g709 (.A(G1399_820_gat), .B(G2213_268_gat), .Y(G1677_909_gat) );
AND2XL U_g710 (.A(G1399_820_gat), .B(G2213_268_gat), .Y(G1929_910_gat) );
AND2XL U_g711 (.A(G1399_820_ngat), .B(G2213_268_ngat), .Y(G5581_911_gat) );
AND2XL U_g712 (.A(G1383_815_gat), .B(G4686_770_gat), .Y(G3015_912_gat) );
BUFX20 U_g713 (.A(G4686_770_gat), .Y(G7463_913_gat) );
BUFX20 U_g714 (.A(G4686_770_gat), .Y(G6431_914_gat) );
INVXL U_g715 (.A(G7466_771_gat), .Y(G7470_915_gat) );
INVXL U_g716 (.A(G6711_772_gat), .Y(G6717_916_gat) );
BUFX20 U_g717 (.A(G1007_773_gat), .Y(G5242_917_gat) );
BUFX20 U_g718 (.A(G1007_773_gat), .Y(G5234_918_gat) );
BUFX20 U_g719 (.A(G765_774_gat), .Y(G4962_919_gat) );
BUFX20 U_g720 (.A(G765_774_gat), .Y(G5003_920_gat) );
INVXL U_g721 (.A(G6714_775_gat), .Y(G6718_921_gat) );
OR2XL U_g722 (.A(G886_604_ngat), .B(G885_832_ngat), .Y(G887_922_gat) );
OR2XL U_g723 (.A(G1018_606_ngat), .B(G1017_831_ngat), .Y(G1019_923_gat) );
AND2XL U_g724 (.A(G2950_865_gat), .B(G1488_279_gat), .Y(G802_924_gat) );
AND2XL U_g725 (.A(G2950_865_gat), .B(G1488_279_gat), .Y(G1035_925_gat) );
AND2XL U_g726 (.A(G645_847_gat), .B(G3679_776_gat), .Y(G3183_926_gat) );
BUFX20 U_g727 (.A(G3679_776_gat), .Y(G6703_927_gat) );
BUFX20 U_g728 (.A(G3679_776_gat), .Y(G6519_928_gat) );
AND2XL U_g729 (.A(G2946_858_gat), .B(G1482_281_gat), .Y(G821_929_gat) );
AND2XL U_g730 (.A(G2946_858_gat), .B(G1482_281_gat), .Y(G1050_930_gat) );
AND2XL U_g731 (.A(G641_841_gat), .B(G3676_777_gat), .Y(G3192_931_gat) );
BUFX20 U_g732 (.A(G3676_777_gat), .Y(G6527_932_gat) );
BUFX20 U_g733 (.A(G3676_777_gat), .Y(G6706_933_gat) );
AND2XL U_g734 (.A(G2938_860_gat), .B(G1471_283_gat), .Y(G868_934_gat) );
AND2XL U_g735 (.A(G2938_860_gat), .B(G1471_283_gat), .Y(G1086_935_gat) );
AND2XL U_g736 (.A(G633_843_gat), .B(G3670_778_gat), .Y(G3207_936_gat) );
BUFX20 U_g737 (.A(G3670_778_gat), .Y(G6543_937_gat) );
BUFX20 U_g738 (.A(G3670_778_gat), .Y(G6698_938_gat) );
AND2XL U_g739 (.A(G2933_861_gat), .B(G1464_285_gat), .Y(G877_939_gat) );
AND2XL U_g740 (.A(G2933_861_gat), .B(G1464_285_gat), .Y(G1102_940_gat) );
AND2XL U_g741 (.A(G2933_861_ngat), .B(G1464_285_ngat), .Y(G5011_941_gat) );
AND2XL U_g742 (.A(G629_844_gat), .B(G3667_779_gat), .Y(G3209_942_gat) );
BUFX20 U_g743 (.A(G3667_779_gat), .Y(G6687_943_gat) );
BUFX20 U_g744 (.A(G3667_779_gat), .Y(G6559_944_gat) );
INVXL U_g745 (.A(G6690_780_gat), .Y(G6694_945_gat) );
INVXL U_g746 (.A(G7296_811_gat), .Y(G7300_946_gat) );
BUFX20 U_g747 (.A(G1387_812_gat), .Y(G6418_947_gat) );
BUFX20 U_g748 (.A(G1387_812_gat), .Y(G7304_948_gat) );
BUFX20 U_g749 (.A(G1391_813_gat), .Y(G7301_949_gat) );
BUFX20 U_g750 (.A(G1391_813_gat), .Y(G6410_950_gat) );
BUFX20 U_g751 (.A(G1395_814_gat), .Y(G6402_951_gat) );
BUFX20 U_g752 (.A(G1395_814_gat), .Y(G7312_952_gat) );
BUFX20 U_g753 (.A(G1383_815_gat), .Y(G7293_953_gat) );
BUFX20 U_g754 (.A(G1383_815_gat), .Y(G6434_954_gat) );
INVXL U_g755 (.A(G5318_816_gat), .Y(G5322_955_gat) );
BUFX20 U_g756 (.A(G1406_817_gat), .Y(G5326_956_gat) );
BUFX20 U_g757 (.A(G1406_817_gat), .Y(G5444_957_gat) );
BUFX20 U_g758 (.A(G1406_817_gat), .Y(G5804_958_gat) );
BUFX20 U_g759 (.A(G1412_818_gat), .Y(G5323_959_gat) );
BUFX20 U_g760 (.A(G1412_818_gat), .Y(G5796_960_gat) );
BUFX20 U_g761 (.A(G1412_818_gat), .Y(G5436_961_gat) );
BUFX20 U_g762 (.A(G1418_819_gat), .Y(G5334_962_gat) );
BUFX20 U_g763 (.A(G1418_819_gat), .Y(G5428_963_gat) );
BUFX20 U_g764 (.A(G1418_819_gat), .Y(G5788_964_gat) );
BUFX20 U_g765 (.A(G1399_820_gat), .Y(G5315_965_gat) );
BUFX20 U_g766 (.A(G1399_820_gat), .Y(G5812_966_gat) );
BUFX20 U_g767 (.A(G1399_820_gat), .Y(G5460_967_gat) );
OR2XL U_g768 (.A(G2048_653_gat), .B(G2047_802_gat), .Y(G2069_968_gat) );
OR2XL U_g769 (.A(G2058_654_gat), .B(G2057_786_gat), .Y(G2091_969_gat) );
OR2XL U_g770 (.A(G2060_655_gat), .B(G2059_787_gat), .Y(G2099_970_gat) );
OR2XL U_g771 (.A(G2050_656_gat), .B(G2049_803_gat), .Y(G2073_971_gat) );
OR2XL U_g772 (.A(G2062_657_gat), .B(G2061_788_gat), .Y(G2105_972_gat) );
OR2XL U_g773 (.A(G2052_658_gat), .B(G2051_804_gat), .Y(G2077_973_gat) );
OR2XL U_g774 (.A(G2162_659_gat), .B(G2161_794_gat), .Y(G2198_974_gat) );
OR2XL U_g775 (.A(G2152_660_gat), .B(G2151_809_gat), .Y(G2175_975_gat) );
OR2XL U_g776 (.A(G2146_661_gat), .B(G2145_810_gat), .Y(G2163_976_gat) );
OR2XL U_g777 (.A(G2156_662_gat), .B(G2155_800_gat), .Y(G2179_977_gat) );
OR2XL U_g778 (.A(G2144_663_gat), .B(G2143_806_gat), .Y(G7208_978_gat) );
OR2XL U_g779 (.A(G2154_664_gat), .B(G2153_791_gat), .Y(G6724_979_gat) );
AND2XL U_g780 (.A(G2942_859_gat), .B(G1477_394_gat), .Y(G845_980_gat) );
AND2XL U_g781 (.A(G2942_859_gat), .B(G1477_394_gat), .Y(G1068_981_gat) );
AND2XL U_g782 (.A(G637_842_gat), .B(G3673_821_gat), .Y(G3200_982_gat) );
BUFX20 U_g783 (.A(G3673_821_gat), .Y(G6695_983_gat) );
BUFX20 U_g784 (.A(G3673_821_gat), .Y(G6535_984_gat) );
OR2XL U_g785 (.A(G2046_673_gat), .B(G2045_801_gat), .Y(G2065_985_gat) );
OR2XL U_g786 (.A(G2056_674_gat), .B(G2055_785_gat), .Y(G2085_986_gat) );
OR2XL U_g787 (.A(G2064_675_gat), .B(G2063_789_gat), .Y(G2111_987_gat) );
OR2XL U_g788 (.A(G2054_676_gat), .B(G2053_805_gat), .Y(G2081_988_gat) );
OR2XL U_g789 (.A(G2158_677_gat), .B(G2157_792_gat), .Y(G2186_989_gat) );
OR2XL U_g790 (.A(G2148_678_gat), .B(G2147_807_gat), .Y(G2167_990_gat) );
OR2XL U_g791 (.A(G2160_679_gat), .B(G2159_793_gat), .Y(G2192_991_gat) );
OR2XL U_g792 (.A(G2150_680_gat), .B(G2149_808_gat), .Y(G2171_992_gat) );
OR2XL U_g793 (.A(G4135_688_gat), .B(G4134_747_gat), .Y(G4160_993_gat) );
OR2XL U_g794 (.A(G4138_689_gat), .B(G4137_746_gat), .Y(G4163_994_gat) );
OR2XL U_g795 (.A(G4141_690_gat), .B(G4140_745_gat), .Y(G4166_995_gat) );
OR2XL U_g796 (.A(G4129_691_gat), .B(G4128_749_gat), .Y(G4154_996_gat) );
OR2XL U_g797 (.A(G4126_692_gat), .B(G4125_750_gat), .Y(G4151_997_gat) );
OR2XL U_g798 (.A(G4477_693_gat), .B(G4476_758_gat), .Y(G4493_998_gat) );
OR2XL U_g799 (.A(G4479_694_gat), .B(G4478_757_gat), .Y(G4496_999_gat) );
OR2XL U_g800 (.A(G4475_695_gat), .B(G4474_759_gat), .Y(G4490_1000_gat) );
OR2XL U_g801 (.A(G4481_696_gat), .B(G4480_756_gat), .Y(G4499_1001_gat) );
OR2XL U_g802 (.A(G4473_697_gat), .B(G4472_760_gat), .Y(G7507_1002_gat) );
OR2XL U_g803 (.A(G4471_699_gat), .B(G4470_761_gat), .Y(G7510_1003_gat) );
OR2XL U_g804 (.A(G3800_700_gat), .B(G3799_799_gat), .Y(G3838_1004_gat) );
BUFX20 U_g805 (.A(G3813_822_gat), .Y(G7239_1005_gat) );
BUFX20 U_g806 (.A(G3813_822_gat), .Y(G6442_1006_gat) );
OR2XL U_g807 (.A(G4150_704_gat), .B(G4149_742_gat), .Y(G4175_1007_gat) );
OR2XL U_g808 (.A(G4147_705_gat), .B(G4146_743_gat), .Y(G4172_1008_gat) );
OR2XL U_g809 (.A(G4144_706_gat), .B(G4143_744_gat), .Y(G4169_1009_gat) );
OR2XL U_g810 (.A(G4132_707_gat), .B(G4131_748_gat), .Y(G4157_1010_gat) );
OR2XL U_g811 (.A(G4123_708_gat), .B(G4122_751_gat), .Y(G7554_1011_gat) );
OR2XL U_g812 (.A(G4489_709_gat), .B(G4488_752_gat), .Y(G4511_1012_gat) );
OR2XL U_g813 (.A(G4487_710_gat), .B(G4486_753_gat), .Y(G4508_1013_gat) );
OR2XL U_g814 (.A(G4485_711_gat), .B(G4484_754_gat), .Y(G4505_1014_gat) );
OR2XL U_g815 (.A(G4483_712_gat), .B(G4482_755_gat), .Y(G4502_1015_gat) );
OR2XL U_g816 (.A(G3798_713_gat), .B(G3797_798_gat), .Y(G3833_1016_gat) );
BUFX20 U_g817 (.A(G3810_823_gat), .Y(G6450_1017_gat) );
BUFX20 U_g818 (.A(G3810_823_gat), .Y(G7242_1018_gat) );
BUFX20 U_g819 (.A(G3801_824_gat), .Y(G6466_1019_gat) );
BUFX20 U_g820 (.A(G3801_824_gat), .Y(G7221_1020_gat) );
OR2XL U_g821 (.A(G3792_714_gat), .B(G3791_795_gat), .Y(G3816_1021_gat) );
INVXL U_g822 (.A(G7252_825_gat), .Y(G7256_1022_gat) );
OR2XL U_g823 (.A(G2296_715_gat), .B(G2295_781_gat), .Y(G6768_1023_gat) );
BUFX20 U_g824 (.A(G2305_826_gat), .Y(G7249_1024_gat) );
OR2XL U_g825 (.A(G2298_716_gat), .B(G2297_790_gat), .Y(G2320_1025_gat) );
OR2XL U_g826 (.A(G6557_741_ngat), .B(G6554_396_ngat), .Y(G3210_1026_gat) );
AND2XL U_g827 (.A(G784_559_gat), .B(G765_774_gat), .Y(G913_1027_gat) );
AND2XL U_g828 (.A(G784_559_gat), .B(G765_774_gat), .Y(G907_1028_gat) );
AND2XL U_g829 (.A(G784_559_gat), .B(G765_774_gat), .Y(G915_1029_gat) );
AND2XL U_g830 (.A(G784_559_gat), .B(G765_774_gat), .Y(G916_1030_gat) );
AND2XL U_g831 (.A(G1014_560_gat), .B(G1007_773_gat), .Y(G1116_1031_gat) );
BUFX20 U_g832 (.A(G3804_833_gat), .Y(G6498_1032_gat) );
BUFX20 U_g833 (.A(G3804_833_gat), .Y(G7232_1033_gat) );
OR2XL U_g834 (.A(G3794_724_gat), .B(G3793_796_gat), .Y(G3821_1034_gat) );
OR2XL U_g835 (.A(G3796_725_gat), .B(G3795_797_gat), .Y(G3828_1035_gat) );
BUFX20 U_g836 (.A(G3807_834_gat), .Y(G6458_1036_gat) );
BUFX20 U_g837 (.A(G3807_834_gat), .Y(G7229_1037_gat) );
OR2XL U_g838 (.A(G2300_726_gat), .B(G2299_782_gat), .Y(G2323_1038_gat) );
BUFX20 U_g839 (.A(G2308_835_gat), .Y(G7412_1039_gat) );
BUFX20 U_g840 (.A(G2308_835_gat), .Y(G7260_1040_gat) );
OR2XL U_g841 (.A(G2302_727_gat), .B(G2301_783_gat), .Y(G2329_1041_gat) );
BUFX20 U_g842 (.A(G2312_836_gat), .Y(G7404_1042_gat) );
BUFX20 U_g843 (.A(G2312_836_gat), .Y(G7257_1043_gat) );
OR2XL U_g844 (.A(G2304_728_gat), .B(G2303_784_gat), .Y(G2335_1044_gat) );
BUFX20 U_g845 (.A(G2316_837_gat), .Y(G7396_1045_gat) );
BUFX20 U_g846 (.A(G2316_837_gat), .Y(G7268_1046_gat) );
BUFX20 U_g847 (.A(G3686_838_gat), .Y(G7425_1047_gat) );
BUFX20 U_g848 (.A(G3682_839_gat), .Y(G5929_1048_gat) );
BUFX20 U_g849 (.A(G3682_839_gat), .Y(G6049_1049_gat) );
AND2XL U_g850 (.A(G2305_826_gat), .B(G1535_302_gat), .Y(G3695_1050_gat) );
INVXL U_g851 (.A(G579_840_gat), .Y(G5284_1051_gat) );
BUFX20 U_g852 (.A(G641_841_gat), .Y(G5300_1052_gat) );
BUFX20 U_g853 (.A(G641_841_gat), .Y(G6530_1053_gat) );
BUFX20 U_g854 (.A(G637_842_gat), .Y(G5289_1054_gat) );
BUFX20 U_g855 (.A(G637_842_gat), .Y(G6538_1055_gat) );
BUFX20 U_g856 (.A(G633_843_gat), .Y(G5292_1056_gat) );
BUFX20 U_g857 (.A(G633_843_gat), .Y(G6546_1057_gat) );
BUFX20 U_g858 (.A(G629_844_gat), .Y(G5281_1058_gat) );
BUFX20 U_g859 (.A(G629_844_gat), .Y(G6562_1059_gat) );
INVXL U_g860 (.A(G5305_845_gat), .Y(G5311_1060_gat) );
INVXL U_g861 (.A(G5308_846_gat), .Y(G5312_1061_gat) );
BUFX20 U_g862 (.A(G645_847_gat), .Y(G5297_1062_gat) );
BUFX20 U_g863 (.A(G645_847_gat), .Y(G6522_1063_gat) );
BUFX20 U_g864 (.A(G727_848_gat), .Y(G7327_1064_gat) );
BUFX20 U_g865 (.A(G727_848_gat), .Y(G6370_1065_gat) );
BUFX20 U_g866 (.A(G723_849_gat), .Y(G6378_1066_gat) );
BUFX20 U_g867 (.A(G723_849_gat), .Y(G7330_1067_gat) );
BUFX20 U_g868 (.A(G719_850_gat), .Y(G7317_1068_gat) );
BUFX20 U_g869 (.A(G719_850_gat), .Y(G6386_1069_gat) );
BUFX20 U_g870 (.A(G715_851_gat), .Y(G6426_1070_gat) );
BUFX20 U_g871 (.A(G715_851_gat), .Y(G7320_1071_gat) );
BUFX20 U_g872 (.A(G711_852_gat), .Y(G7309_1072_gat) );
BUFX20 U_g873 (.A(G711_852_gat), .Y(G6394_1073_gat) );
BUFX20 U_g874 (.A(G745_853_gat), .Y(G5339_1074_gat) );
BUFX20 U_g875 (.A(G745_853_gat), .Y(G5764_1075_gat) );
BUFX20 U_g876 (.A(G745_853_gat), .Y(G5412_1076_gat) );
BUFX20 U_g877 (.A(G737_854_gat), .Y(G5452_1077_gat) );
BUFX20 U_g878 (.A(G737_854_gat), .Y(G5772_1078_gat) );
BUFX20 U_g879 (.A(G737_854_gat), .Y(G5342_1079_gat) );
BUFX20 U_g880 (.A(G731_855_gat), .Y(G5331_1080_gat) );
BUFX20 U_g881 (.A(G731_855_gat), .Y(G5780_1081_gat) );
BUFX20 U_g882 (.A(G731_855_gat), .Y(G5420_1082_gat) );
BUFX20 U_g883 (.A(G757_856_gat), .Y(G5349_1083_gat) );
BUFX20 U_g884 (.A(G757_856_gat), .Y(G5396_1084_gat) );
BUFX20 U_g885 (.A(G757_856_gat), .Y(G5748_1085_gat) );
BUFX20 U_g886 (.A(G751_857_gat), .Y(G5756_1086_gat) );
BUFX20 U_g887 (.A(G751_857_gat), .Y(G5404_1087_gat) );
BUFX20 U_g888 (.A(G751_857_gat), .Y(G5352_1088_gat) );
BUFX20 U_g889 (.A(G2946_858_gat), .Y(G5202_1089_gat) );
BUFX20 U_g890 (.A(G2946_858_gat), .Y(G4892_1090_gat) );
BUFX20 U_g891 (.A(G2946_858_gat), .Y(G5266_1091_gat) );
BUFX20 U_g892 (.A(G2942_859_gat), .Y(G5255_1092_gat) );
BUFX20 U_g893 (.A(G2942_859_gat), .Y(G4900_1093_gat) );
BUFX20 U_g894 (.A(G2942_859_gat), .Y(G5210_1094_gat) );
BUFX20 U_g895 (.A(G2938_860_gat), .Y(G5218_1095_gat) );
BUFX20 U_g896 (.A(G2938_860_gat), .Y(G4908_1096_gat) );
BUFX20 U_g897 (.A(G2938_860_gat), .Y(G5258_1097_gat) );
BUFX20 U_g898 (.A(G2933_861_gat), .Y(G5247_1098_gat) );
BUFX20 U_g899 (.A(G2933_861_gat), .Y(G4924_1099_gat) );
BUFX20 U_g900 (.A(G2933_861_gat), .Y(G5226_1100_gat) );
INVXL U_g901 (.A(G4525_862_gat), .Y(G5250_1101_gat) );
INVXL U_g902 (.A(G5271_863_gat), .Y(G5277_1102_gat) );
INVXL U_g903 (.A(G5274_864_gat), .Y(G5278_1103_gat) );
BUFX20 U_g904 (.A(G2950_865_gat), .Y(G5263_1104_gat) );
BUFX20 U_g905 (.A(G2950_865_gat), .Y(G4884_1105_gat) );
BUFX20 U_g906 (.A(G2950_865_gat), .Y(G5194_1106_gat) );
AND2XL U_g907 (.A(G3838_1004_gat), .B(G4439_209_gat), .Y(G3292_1107_gat) );
AND2XL U_g908 (.A(G3838_1004_gat), .B(G4439_209_gat), .Y(G3853_1108_gat) );
AND2XL U_g909 (.A(G3833_1016_gat), .B(G4434_211_gat), .Y(G3308_1109_gat) );
AND2XL U_g910 (.A(G3833_1016_gat), .B(G4434_211_gat), .Y(G3868_1110_gat) );
AND2XL U_g911 (.A(G3828_1035_gat), .B(G4429_213_gat), .Y(G3327_1111_gat) );
AND2XL U_g912 (.A(G3828_1035_gat), .B(G4429_213_gat), .Y(G3885_1112_gat) );
AND2XL U_g913 (.A(G4422_215_gat), .B(G3821_1034_gat), .Y(G3335_1113_gat) );
AND2XL U_g914 (.A(G3821_1034_gat), .B(G4422_215_gat), .Y(G3891_1114_gat) );
AND2XL U_g915 (.A(G3821_1034_ngat), .B(G4422_215_ngat), .Y(G6925_1115_gat) );
AND2XL U_g916 (.A(G4422_215_ngat), .B(G3821_1034_ngat), .Y(G6671_1116_gat) );
AND2XL U_g917 (.A(G3816_1021_gat), .B(G4417_217_gat), .Y(G3362_1117_gat) );
AND2XL U_g918 (.A(G3816_1021_gat), .B(G4417_217_gat), .Y(G3908_1118_gat) );
AND2XL U_g919 (.A(G2198_974_gat), .B(G4412_219_gat), .Y(G3376_1119_gat) );
AND2XL U_g920 (.A(G2198_974_gat), .B(G4412_219_gat), .Y(G3926_1120_gat) );
AND2XL U_g921 (.A(G2192_991_gat), .B(G4407_221_gat), .Y(G3393_1121_gat) );
AND2XL U_g922 (.A(G2192_991_gat), .B(G4407_221_gat), .Y(G3949_1122_gat) );
AND2XL U_g923 (.A(G2186_989_gat), .B(G4402_223_gat), .Y(G3410_1123_gat) );
AND2XL U_g924 (.A(G2186_989_gat), .B(G4402_223_gat), .Y(G3971_1124_gat) );
AND2XL U_g925 (.A(G2179_977_gat), .B(G4396_225_gat), .Y(G3425_1125_gat) );
AND2XL U_g926 (.A(G2179_977_gat), .B(G4396_225_gat), .Y(G3979_1126_gat) );
AND2XL U_g927 (.A(G2179_977_ngat), .B(G4396_225_ngat), .Y(G7041_1127_gat) );
AND2XL U_g928 (.A(G2111_987_gat), .B(G3751_229_gat), .Y(G2351_1128_gat) );
AND2XL U_g929 (.A(G2111_987_gat), .B(G3751_229_gat), .Y(G2597_1129_gat) );
AND2XL U_g930 (.A(G2105_972_gat), .B(G3745_231_gat), .Y(G2366_1130_gat) );
AND2XL U_g931 (.A(G2105_972_gat), .B(G3745_231_gat), .Y(G2612_1131_gat) );
AND2XL U_g932 (.A(G2099_970_gat), .B(G3739_233_gat), .Y(G2384_1132_gat) );
AND2XL U_g933 (.A(G2099_970_gat), .B(G3739_233_gat), .Y(G2629_1133_gat) );
AND2XL U_g934 (.A(G3731_235_gat), .B(G2091_969_gat), .Y(G2391_1134_gat) );
AND2XL U_g935 (.A(G2091_969_gat), .B(G3731_235_gat), .Y(G2635_1135_gat) );
AND2XL U_g936 (.A(G2091_969_ngat), .B(G3731_235_ngat), .Y(G6057_1136_gat) );
AND2XL U_g937 (.A(G3731_235_ngat), .B(G2091_969_ngat), .Y(G5969_1137_gat) );
AND2XL U_g938 (.A(G2085_986_gat), .B(G3725_237_gat), .Y(G2417_1138_gat) );
AND2XL U_g939 (.A(G2085_986_gat), .B(G3725_237_gat), .Y(G2652_1139_gat) );
AND2XL U_g940 (.A(G2335_1044_gat), .B(G3719_239_gat), .Y(G2431_1140_gat) );
AND2XL U_g941 (.A(G2335_1044_gat), .B(G3719_239_gat), .Y(G2670_1141_gat) );
AND2XL U_g942 (.A(G2329_1041_gat), .B(G3713_241_gat), .Y(G2448_1142_gat) );
AND2XL U_g943 (.A(G2329_1041_gat), .B(G3713_241_gat), .Y(G2693_1143_gat) );
AND2XL U_g944 (.A(G2323_1038_gat), .B(G3707_243_gat), .Y(G2465_1144_gat) );
AND2XL U_g945 (.A(G2323_1038_gat), .B(G3707_243_gat), .Y(G2715_1145_gat) );
INVXL U_g946 (.A(G7497_868_gat), .Y(G7503_1146_gat) );
INVXL U_g947 (.A(G6367_869_gat), .Y(G6373_1147_gat) );
OR2XL U_g948 (.A(G5399_466_ngat), .B(G5396_1084_ngat), .Y(G1544_1148_gat) );
OR2XL U_g949 (.A(G5751_467_ngat), .B(G5748_1085_ngat), .Y(G1793_1149_gat) );
INVXL U_g950 (.A(G7500_873_gat), .Y(G7504_1150_gat) );
INVXL U_g951 (.A(G6375_874_gat), .Y(G6381_1151_gat) );
OR2XL U_g952 (.A(G5759_469_ngat), .B(G5756_1086_ngat), .Y(G1803_1152_gat) );
OR2XL U_g953 (.A(G5407_470_ngat), .B(G5404_1087_ngat), .Y(G1554_1153_gat) );
INVXL U_g954 (.A(G6383_880_gat), .Y(G6389_1154_gat) );
INVXL U_g955 (.A(G7487_881_gat), .Y(G7493_1155_gat) );
OR2XL U_g956 (.A(G5415_472_ngat), .B(G5412_1076_ngat), .Y(G1571_1156_gat) );
OR2XL U_g957 (.A(G5767_473_ngat), .B(G5764_1075_ngat), .Y(G1820_1157_gat) );
BUFX20 U_g958 (.A(G1590_882_gat), .Y(G5523_1158_gat) );
BUFX20 U_g959 (.A(G1841_883_gat), .Y(G5857_1159_gat) );
OR2XL U_g960 (.A(G5775_474_ngat), .B(G5772_1078_ngat), .Y(G1848_1160_gat) );
INVXL U_g961 (.A(G5849_884_gat), .Y(G5855_1161_gat) );
INVXL U_g962 (.A(G5465_885_gat), .Y(G5471_1162_gat) );
OR2XL U_g963 (.A(G5455_475_ngat), .B(G5452_1077_ngat), .Y(G1685_1163_gat) );
INVXL U_g964 (.A(G7490_887_gat), .Y(G7494_1164_gat) );
INVXL U_g965 (.A(G6423_888_gat), .Y(G6429_1165_gat) );
INVXL U_g966 (.A(G7479_890_gat), .Y(G7485_1166_gat) );
INVXL U_g967 (.A(G6391_891_gat), .Y(G6397_1167_gat) );
OR2XL U_g968 (.A(G5423_478_ngat), .B(G5420_1082_ngat), .Y(G1596_1168_gat) );
OR2XL U_g969 (.A(G5783_479_ngat), .B(G5780_1081_ngat), .Y(G1857_1169_gat) );
OR2XL U_g970 (.A(G5791_480_ngat), .B(G5788_964_ngat), .Y(G1867_1170_gat) );
OR2XL U_g971 (.A(G5431_481_ngat), .B(G5428_963_ngat), .Y(G1607_1171_gat) );
INVXL U_g972 (.A(G6399_897_gat), .Y(G6405_1172_gat) );
INVXL U_g973 (.A(G7482_898_gat), .Y(G7486_1173_gat) );
INVXL U_g974 (.A(G7471_902_gat), .Y(G7477_1174_gat) );
INVXL U_g975 (.A(G6407_903_gat), .Y(G6413_1175_gat) );
OR2XL U_g976 (.A(G5439_484_ngat), .B(G5436_961_ngat), .Y(G1628_1176_gat) );
OR2XL U_g977 (.A(G5799_485_ngat), .B(G5796_960_ngat), .Y(G1883_1177_gat) );
OR2XL U_g978 (.A(G5807_486_ngat), .B(G5804_958_ngat), .Y(G1901_1178_gat) );
OR2XL U_g979 (.A(G5447_487_ngat), .B(G5444_957_ngat), .Y(G1653_1179_gat) );
INVXL U_g980 (.A(G6415_907_gat), .Y(G6421_1180_gat) );
INVXL U_g981 (.A(G7474_908_gat), .Y(G7478_1181_gat) );
BUFX20 U_g982 (.A(G1677_909_gat), .Y(G5669_1182_gat) );
INVXL U_g983 (.A(G5581_911_gat), .Y(G5587_1183_gat) );
OR2XL U_g984 (.A(G5463_489_ngat), .B(G5460_967_ngat), .Y(G1693_1184_gat) );
OR2XL U_g985 (.A(G7470_915_ngat), .B(G7463_913_ngat), .Y(G4530_1185_gat) );
INVXL U_g986 (.A(G7463_913_gat), .Y(G7469_1186_gat) );
INVXL U_g987 (.A(G6431_914_gat), .Y(G6437_1187_gat) );
OR2XL U_g988 (.A(G5815_491_ngat), .B(G5812_966_ngat), .Y(G1919_1188_gat) );
OR2XL U_g989 (.A(G6718_921_ngat), .B(G6711_772_ngat), .Y(G6720_1189_gat) );
OR2XL U_g990 (.A(G916_1030_gat), .B(G777_370_gat), .Y(G917_1190_gat) );
AND2XL U_g991 (.A(G915_1029_ngat), .B(G777_370_ngat), .Y(G4983_1191_gat) );
OR2XL U_g992 (.A(G907_1028_gat), .B(G777_370_gat), .Y(G908_1192_gat) );
OR2XL U_g993 (.A(G1116_1031_gat), .B(G1115_371_gat), .Y(G1117_1193_gat) );
INVXL U_g994 (.A(G5242_917_gat), .Y(G5246_1194_gat) );
INVXL U_g995 (.A(G5234_918_gat), .Y(G5238_1195_gat) );
AND2XL U_g996 (.A(G1007_773_gat), .B(G1019_923_gat), .Y(G1108_1196_gat) );
AND2XL U_g997 (.A(G765_774_gat), .B(G887_922_gat), .Y(G953_1197_gat) );
INVXL U_g998 (.A(G4962_919_gat), .Y(G4966_1198_gat) );
AND2XL U_g999 (.A(G765_774_gat), .B(G887_922_gat), .Y(G902_1199_gat) );
AND2XL U_g1000 (.A(G765_774_gat), .B(G887_922_gat), .Y(G914_1200_gat) );
INVXL U_g1001 (.A(G5003_920_gat), .Y(G5007_1201_gat) );
OR2XL U_g1002 (.A(G6717_916_ngat), .B(G6714_775_ngat), .Y(G6719_1202_gat) );
BUFX20 U_g1003 (.A(G887_922_gat), .Y(G4993_1203_gat) );
BUFX20 U_g1004 (.A(G887_922_gat), .Y(G4952_1204_gat) );
INVXL U_g1005 (.A(G1019_923_gat), .Y(G1023_1205_gat) );
INVXL U_g1006 (.A(G6703_927_gat), .Y(G6709_1206_gat) );
INVXL U_g1007 (.A(G6519_928_gat), .Y(G6525_1207_gat) );
OR2XL U_g1008 (.A(G4887_500_ngat), .B(G4884_1105_ngat), .Y(G790_1208_gat) );
OR2XL U_g1009 (.A(G5197_501_ngat), .B(G5194_1106_ngat), .Y(G1024_1209_gat) );
OR2XL U_g1010 (.A(G5205_502_ngat), .B(G5202_1089_ngat), .Y(G1036_1210_gat) );
OR2XL U_g1011 (.A(G4895_503_ngat), .B(G4892_1090_ngat), .Y(G803_1211_gat) );
INVXL U_g1012 (.A(G6527_932_gat), .Y(G6533_1212_gat) );
INVXL U_g1013 (.A(G6706_933_gat), .Y(G6710_1213_gat) );
OR2XL U_g1014 (.A(G5221_505_ngat), .B(G5218_1095_ngat), .Y(G1072_1214_gat) );
INVXL U_g1015 (.A(G6543_937_gat), .Y(G6549_1215_gat) );
INVXL U_g1016 (.A(G6698_938_gat), .Y(G6702_1216_gat) );
OR2XL U_g1017 (.A(G4911_507_ngat), .B(G4908_1096_ngat), .Y(G851_1217_gat) );
BUFX20 U_g1018 (.A(G877_939_gat), .Y(G5099_1218_gat) );
INVXL U_g1019 (.A(G5011_941_gat), .Y(G5017_1219_gat) );
OR2XL U_g1020 (.A(G4927_508_ngat), .B(G4924_1099_ngat), .Y(G893_1220_gat) );
OR2XL U_g1021 (.A(G6694_945_ngat), .B(G6687_943_ngat), .Y(G3503_1221_gat) );
INVXL U_g1022 (.A(G6687_943_gat), .Y(G6693_1222_gat) );
INVXL U_g1023 (.A(G6559_944_gat), .Y(G6565_1223_gat) );
OR2XL U_g1024 (.A(G5229_510_ngat), .B(G5226_1100_ngat), .Y(G1091_1224_gat) );
OR2XL U_g1025 (.A(G7300_946_ngat), .B(G7293_953_ngat), .Y(G4225_1225_gat) );
INVXL U_g1026 (.A(G6418_947_gat), .Y(G6422_1226_gat) );
INVXL U_g1027 (.A(G7304_948_gat), .Y(G7308_1227_gat) );
INVXL U_g1028 (.A(G7301_949_gat), .Y(G7307_1228_gat) );
INVXL U_g1029 (.A(G6410_950_gat), .Y(G6414_1229_gat) );
INVXL U_g1030 (.A(G6402_951_gat), .Y(G6406_1230_gat) );
INVXL U_g1031 (.A(G7312_952_gat), .Y(G7316_1231_gat) );
INVXL U_g1032 (.A(G7293_953_gat), .Y(G7299_1232_gat) );
INVXL U_g1033 (.A(G6434_954_gat), .Y(G6438_1233_gat) );
OR2XL U_g1034 (.A(G5322_955_ngat), .B(G5315_965_ngat), .Y(G1262_1234_gat) );
INVXL U_g1035 (.A(G5326_956_gat), .Y(G5330_1235_gat) );
INVXL U_g1036 (.A(G5444_957_gat), .Y(G5448_1236_gat) );
INVXL U_g1037 (.A(G5804_958_gat), .Y(G5808_1237_gat) );
INVXL U_g1038 (.A(G5323_959_gat), .Y(G5329_1238_gat) );
INVXL U_g1039 (.A(G5796_960_gat), .Y(G5800_1239_gat) );
INVXL U_g1040 (.A(G5436_961_gat), .Y(G5440_1240_gat) );
INVXL U_g1041 (.A(G5334_962_gat), .Y(G5338_1241_gat) );
INVXL U_g1042 (.A(G5428_963_gat), .Y(G5432_1242_gat) );
INVXL U_g1043 (.A(G5788_964_gat), .Y(G5792_1243_gat) );
INVXL U_g1044 (.A(G5315_965_gat), .Y(G5321_1244_gat) );
INVXL U_g1045 (.A(G5812_966_gat), .Y(G5816_1245_gat) );
INVXL U_g1046 (.A(G5460_967_gat), .Y(G5464_1246_gat) );
BUFX20 U_g1047 (.A(G2069_968_gat), .Y(G7276_1247_gat) );
AND2XL U_g1048 (.A(G2069_968_gat), .B(G4502_1015_gat), .Y(G4314_1248_gat) );
BUFX20 U_g1049 (.A(G2069_968_gat), .Y(G7420_1249_gat) );
BUFX20 U_g1050 (.A(G2091_969_gat), .Y(G5892_1250_gat) );
BUFX20 U_g1051 (.A(G2091_969_gat), .Y(G6044_1251_gat) );
BUFX20 U_g1052 (.A(G2091_969_gat), .Y(G6792_1252_gat) );
BUFX20 U_g1053 (.A(G2099_970_gat), .Y(G6789_1253_gat) );
BUFX20 U_g1054 (.A(G2099_970_gat), .Y(G6004_1254_gat) );
BUFX20 U_g1055 (.A(G2099_970_gat), .Y(G5884_1255_gat) );
AND2XL U_g1056 (.A(G2073_971_gat), .B(G4505_1014_gat), .Y(G4312_1256_gat) );
BUFX20 U_g1057 (.A(G2073_971_gat), .Y(G7380_1257_gat) );
BUFX20 U_g1058 (.A(G2073_971_gat), .Y(G7273_1258_gat) );
BUFX20 U_g1059 (.A(G2105_972_gat), .Y(G5876_1259_gat) );
BUFX20 U_g1060 (.A(G2105_972_gat), .Y(G5996_1260_gat) );
BUFX20 U_g1061 (.A(G2105_972_gat), .Y(G6802_1261_gat) );
AND2XL U_g1062 (.A(G2077_973_gat), .B(G4508_1013_gat), .Y(G4305_1262_gat) );
BUFX20 U_g1063 (.A(G2077_973_gat), .Y(G7372_1263_gat) );
BUFX20 U_g1064 (.A(G2077_973_gat), .Y(G7286_1264_gat) );
BUFX20 U_g1065 (.A(G2198_974_gat), .Y(G6740_1265_gat) );
BUFX20 U_g1066 (.A(G2198_974_gat), .Y(G6610_1266_gat) );
BUFX20 U_g1067 (.A(G2198_974_gat), .Y(G6888_1267_gat) );
AND2XL U_g1068 (.A(G2175_975_gat), .B(G4160_993_gat), .Y(G3099_1268_gat) );
BUFX20 U_g1069 (.A(G2175_975_gat), .Y(G6474_1269_gat) );
BUFX20 U_g1070 (.A(G2175_975_gat), .Y(G7224_1270_gat) );
AND2XL U_g1071 (.A(G2163_976_gat), .B(G4151_997_gat), .Y(G3116_1271_gat) );
BUFX20 U_g1072 (.A(G2163_976_gat), .Y(G6506_1272_gat) );
BUFX20 U_g1073 (.A(G2163_976_gat), .Y(G7205_1273_gat) );
BUFX20 U_g1074 (.A(G2179_977_gat), .Y(G6721_1274_gat) );
BUFX20 U_g1075 (.A(G2179_977_gat), .Y(G6634_1275_gat) );
BUFX20 U_g1076 (.A(G2179_977_gat), .Y(G6920_1276_gat) );
INVXL U_g1077 (.A(G7208_978_gat), .Y(G7212_1277_gat) );
INVXL U_g1078 (.A(G6724_979_gat), .Y(G6728_1278_gat) );
OR2XL U_g1079 (.A(G4903_671_ngat), .B(G4900_1093_ngat), .Y(G825_1279_gat) );
OR2XL U_g1080 (.A(G5213_672_ngat), .B(G5210_1094_ngat), .Y(G1053_1280_gat) );
INVXL U_g1081 (.A(G6695_983_gat), .Y(G6701_1281_gat) );
INVXL U_g1082 (.A(G6535_984_gat), .Y(G6541_1282_gat) );
BUFX20 U_g1083 (.A(G2065_985_gat), .Y(G7388_1283_gat) );
AND2XL U_g1084 (.A(G2065_985_gat), .B(G4499_1001_gat), .Y(G4324_1284_gat) );
BUFX20 U_g1085 (.A(G2065_985_gat), .Y(G7265_1285_gat) );
BUFX20 U_g1086 (.A(G2085_986_gat), .Y(G6781_1286_gat) );
BUFX20 U_g1087 (.A(G2085_986_gat), .Y(G6012_1287_gat) );
BUFX20 U_g1088 (.A(G2085_986_gat), .Y(G5900_1288_gat) );
BUFX20 U_g1089 (.A(G2111_987_gat), .Y(G6799_1289_gat) );
BUFX20 U_g1090 (.A(G2111_987_gat), .Y(G5988_1290_gat) );
BUFX20 U_g1091 (.A(G2111_987_gat), .Y(G5868_1291_gat) );
BUFX20 U_g1092 (.A(G2081_988_gat), .Y(G7364_1292_gat) );
AND2XL U_g1093 (.A(G2081_988_gat), .B(G4511_1012_gat), .Y(G4297_1293_gat) );
BUFX20 U_g1094 (.A(G2081_988_gat), .Y(G7283_1294_gat) );
BUFX20 U_g1095 (.A(G2186_989_gat), .Y(G6732_1295_gat) );
BUFX20 U_g1096 (.A(G2186_989_gat), .Y(G6904_1296_gat) );
BUFX20 U_g1097 (.A(G2186_989_gat), .Y(G6626_1297_gat) );
AND2XL U_g1098 (.A(G2167_990_gat), .B(G4154_996_gat), .Y(G3114_1298_gat) );
BUFX20 U_g1099 (.A(G2167_990_gat), .Y(G6490_1299_gat) );
BUFX20 U_g1100 (.A(G2167_990_gat), .Y(G7216_1300_gat) );
BUFX20 U_g1101 (.A(G2192_991_gat), .Y(G6729_1301_gat) );
BUFX20 U_g1102 (.A(G2192_991_gat), .Y(G6896_1302_gat) );
BUFX20 U_g1103 (.A(G2192_991_gat), .Y(G6618_1303_gat) );
BUFX20 U_g1104 (.A(G2171_992_gat), .Y(G6482_1304_gat) );
AND2XL U_g1105 (.A(G2171_992_gat), .B(G4157_1010_gat), .Y(G3107_1305_gat) );
BUFX20 U_g1106 (.A(G2171_992_gat), .Y(G7213_1306_gat) );
BUFX20 U_g1107 (.A(G4160_993_gat), .Y(G6471_1307_gat) );
BUFX20 U_g1108 (.A(G4160_993_gat), .Y(G7570_1308_gat) );
BUFX20 U_g1109 (.A(G4163_994_gat), .Y(G6463_1309_gat) );
BUFX20 U_g1110 (.A(G4163_994_gat), .Y(G7567_1310_gat) );
BUFX20 U_g1111 (.A(G4166_995_gat), .Y(G6495_1311_gat) );
BUFX20 U_g1112 (.A(G4166_995_gat), .Y(G7578_1312_gat) );
BUFX20 U_g1113 (.A(G4154_996_gat), .Y(G6487_1313_gat) );
BUFX20 U_g1114 (.A(G4154_996_gat), .Y(G7562_1314_gat) );
BUFX20 U_g1115 (.A(G4151_997_gat), .Y(G6503_1315_gat) );
BUFX20 U_g1116 (.A(G4151_997_gat), .Y(G7551_1316_gat) );
BUFX20 U_g1117 (.A(G4493_998_gat), .Y(G7515_1317_gat) );
BUFX20 U_g1118 (.A(G4493_998_gat), .Y(G7401_1318_gat) );
BUFX20 U_g1119 (.A(G4496_999_gat), .Y(G7393_1319_gat) );
BUFX20 U_g1120 (.A(G4496_999_gat), .Y(G7526_1320_gat) );
BUFX20 U_g1121 (.A(G4490_1000_gat), .Y(G7409_1321_gat) );
BUFX20 U_g1122 (.A(G4490_1000_gat), .Y(G7518_1322_gat) );
BUFX20 U_g1123 (.A(G4499_1001_gat), .Y(G7523_1323_gat) );
BUFX20 U_g1124 (.A(G4499_1001_gat), .Y(G7385_1324_gat) );
INVXL U_g1125 (.A(G7507_1002_gat), .Y(G7513_1325_gat) );
INVXL U_g1126 (.A(G7510_1003_gat), .Y(G7514_1326_gat) );
BUFX20 U_g1127 (.A(G3838_1004_gat), .Y(G6856_1327_gat) );
BUFX20 U_g1128 (.A(G3838_1004_gat), .Y(G6755_1328_gat) );
BUFX20 U_g1129 (.A(G3838_1004_gat), .Y(G6570_1329_gat) );
AND2XL U_g1130 (.A(G3813_822_gat), .B(G4175_1007_gat), .Y(G3059_1330_gat) );
INVXL U_g1131 (.A(G7239_1005_gat), .Y(G7245_1331_gat) );
INVXL U_g1132 (.A(G6442_1006_gat), .Y(G6446_1332_gat) );
BUFX20 U_g1133 (.A(G4175_1007_gat), .Y(G6439_1333_gat) );
BUFX20 U_g1134 (.A(G4175_1007_gat), .Y(G7585_1334_gat) );
BUFX20 U_g1135 (.A(G4172_1008_gat), .Y(G6447_1335_gat) );
BUFX20 U_g1136 (.A(G4172_1008_gat), .Y(G7588_1336_gat) );
BUFX20 U_g1137 (.A(G4169_1009_gat), .Y(G6455_1337_gat) );
BUFX20 U_g1138 (.A(G4169_1009_gat), .Y(G7575_1338_gat) );
BUFX20 U_g1139 (.A(G4157_1010_gat), .Y(G6479_1339_gat) );
BUFX20 U_g1140 (.A(G4157_1010_gat), .Y(G7559_1340_gat) );
INVXL U_g1141 (.A(G7554_1011_gat), .Y(G7558_1341_gat) );
BUFX20 U_g1142 (.A(G4511_1012_gat), .Y(G7541_1342_gat) );
BUFX20 U_g1143 (.A(G4511_1012_gat), .Y(G7361_1343_gat) );
BUFX20 U_g1144 (.A(G4508_1013_gat), .Y(G7369_1344_gat) );
BUFX20 U_g1145 (.A(G4508_1013_gat), .Y(G7544_1345_gat) );
BUFX20 U_g1146 (.A(G4505_1014_gat), .Y(G7531_1346_gat) );
BUFX20 U_g1147 (.A(G4505_1014_gat), .Y(G7377_1347_gat) );
BUFX20 U_g1148 (.A(G4502_1015_gat), .Y(G7534_1348_gat) );
BUFX20 U_g1149 (.A(G4502_1015_gat), .Y(G7417_1349_gat) );
BUFX20 U_g1150 (.A(G3833_1016_gat), .Y(G6578_1350_gat) );
BUFX20 U_g1151 (.A(G3833_1016_gat), .Y(G6758_1351_gat) );
BUFX20 U_g1152 (.A(G3833_1016_gat), .Y(G6864_1352_gat) );
AND2XL U_g1153 (.A(G3810_823_gat), .B(G4172_1008_gat), .Y(G3068_1353_gat) );
INVXL U_g1154 (.A(G6450_1017_gat), .Y(G6454_1354_gat) );
INVXL U_g1155 (.A(G7242_1018_gat), .Y(G7246_1355_gat) );
AND2XL U_g1156 (.A(G3801_824_gat), .B(G4163_994_gat), .Y(G3090_1356_gat) );
INVXL U_g1157 (.A(G6466_1019_gat), .Y(G6470_1357_gat) );
INVXL U_g1158 (.A(G7221_1020_gat), .Y(G7227_1358_gat) );
BUFX20 U_g1159 (.A(G3816_1021_gat), .Y(G6602_1359_gat) );
BUFX20 U_g1160 (.A(G3816_1021_gat), .Y(G6737_1360_gat) );
BUFX20 U_g1161 (.A(G3816_1021_gat), .Y(G6880_1361_gat) );
OR2XL U_g1162 (.A(G7256_1022_ngat), .B(G7249_1024_ngat), .Y(G4202_1362_gat) );
INVXL U_g1163 (.A(G6768_1023_gat), .Y(G6772_1363_gat) );
INVXL U_g1164 (.A(G7249_1024_gat), .Y(G7255_1364_gat) );
BUFX20 U_g1165 (.A(G2320_1025_gat), .Y(G6765_1365_gat) );
AND2XL U_g1166 (.A(G3173_717_gat), .B(G3170_866_gat), .Y(G3222_1366_gat) );
OR2XL U_g1167 (.A(G3211_827_ngat), .B(G3210_1026_ngat), .Y(G3212_1367_gat) );
OR2XL U_g1168 (.A(G5245_830_ngat), .B(G5242_917_ngat), .Y(G1156_1368_gat) );
OR2XL U_g1169 (.A(G5237_720_ngat), .B(G5234_918_ngat), .Y(G1152_1369_gat) );
AND2XL U_g1170 (.A(G3804_833_gat), .B(G4166_995_gat), .Y(G3079_1370_gat) );
INVXL U_g1171 (.A(G6498_1032_gat), .Y(G6502_1371_gat) );
INVXL U_g1172 (.A(G7232_1033_gat), .Y(G7236_1372_gat) );
BUFX20 U_g1173 (.A(G3821_1034_gat), .Y(G6748_1373_gat) );
BUFX20 U_g1174 (.A(G3821_1034_gat), .Y(G6912_1374_gat) );
BUFX20 U_g1175 (.A(G3821_1034_gat), .Y(G6594_1375_gat) );
BUFX20 U_g1176 (.A(G3828_1035_gat), .Y(G6745_1376_gat) );
BUFX20 U_g1177 (.A(G3828_1035_gat), .Y(G6872_1377_gat) );
BUFX20 U_g1178 (.A(G3828_1035_gat), .Y(G6586_1378_gat) );
AND2XL U_g1179 (.A(G3807_834_gat), .B(G4169_1009_gat), .Y(G3076_1379_gat) );
INVXL U_g1180 (.A(G6458_1036_gat), .Y(G6462_1380_gat) );
INVXL U_g1181 (.A(G7229_1037_gat), .Y(G7235_1381_gat) );
BUFX20 U_g1182 (.A(G2323_1038_gat), .Y(G5924_1382_gat) );
BUFX20 U_g1183 (.A(G2323_1038_gat), .Y(G6036_1383_gat) );
BUFX20 U_g1184 (.A(G2323_1038_gat), .Y(G6776_1384_gat) );
AND2XL U_g1185 (.A(G2308_835_gat), .B(G4490_1000_gat), .Y(G4348_1385_gat) );
INVXL U_g1186 (.A(G7412_1039_gat), .Y(G7416_1386_gat) );
INVXL U_g1187 (.A(G7260_1040_gat), .Y(G7264_1387_gat) );
BUFX20 U_g1188 (.A(G2329_1041_gat), .Y(G6773_1388_gat) );
BUFX20 U_g1189 (.A(G2329_1041_gat), .Y(G6028_1389_gat) );
BUFX20 U_g1190 (.A(G2329_1041_gat), .Y(G5916_1390_gat) );
INVXL U_g1191 (.A(G7404_1042_gat), .Y(G7408_1391_gat) );
AND2XL U_g1192 (.A(G2312_836_gat), .B(G4493_998_gat), .Y(G4341_1392_gat) );
INVXL U_g1193 (.A(G7257_1043_gat), .Y(G7263_1393_gat) );
BUFX20 U_g1194 (.A(G2335_1044_gat), .Y(G5908_1394_gat) );
BUFX20 U_g1195 (.A(G2335_1044_gat), .Y(G6020_1395_gat) );
BUFX20 U_g1196 (.A(G2335_1044_gat), .Y(G6784_1396_gat) );
AND2XL U_g1197 (.A(G2316_837_gat), .B(G4496_999_gat), .Y(G4333_1397_gat) );
INVXL U_g1198 (.A(G7396_1045_gat), .Y(G7400_1398_gat) );
INVXL U_g1199 (.A(G7268_1046_gat), .Y(G7272_1399_gat) );
AND2XL U_g1200 (.A(G3695_1050_gat), .B(G3686_838_gat), .Y(G4349_1400_gat) );
INVXL U_g1201 (.A(G7425_1047_gat), .Y(G7431_1401_gat) );
INVXL U_g1202 (.A(G5929_1048_gat), .Y(G5935_1402_gat) );
INVXL U_g1203 (.A(G6049_1049_gat), .Y(G6055_1403_gat) );
BUFX20 U_g1204 (.A(G3695_1050_gat), .Y(G7428_1404_gat) );
AND2XL U_g1205 (.A(G1535_302_gat), .B(G2320_1025_gat), .Y(G4389_1405_gat) );
INVXL U_g1206 (.A(G5284_1051_gat), .Y(G5288_1406_gat) );
INVXL U_g1207 (.A(G5300_1052_gat), .Y(G5304_1407_gat) );
INVXL U_g1208 (.A(G6530_1053_gat), .Y(G6534_1408_gat) );
INVXL U_g1209 (.A(G5289_1054_gat), .Y(G5295_1409_gat) );
INVXL U_g1210 (.A(G6538_1055_gat), .Y(G6542_1410_gat) );
INVXL U_g1211 (.A(G5292_1056_gat), .Y(G5296_1411_gat) );
INVXL U_g1212 (.A(G6546_1057_gat), .Y(G6550_1412_gat) );
INVXL U_g1213 (.A(G5281_1058_gat), .Y(G5287_1413_gat) );
INVXL U_g1214 (.A(G6562_1059_gat), .Y(G6566_1414_gat) );
OR2XL U_g1215 (.A(G5312_1061_ngat), .B(G5305_845_ngat), .Y(G5314_1415_gat) );
OR2XL U_g1216 (.A(G5311_1060_ngat), .B(G5308_846_ngat), .Y(G5313_1416_gat) );
INVXL U_g1217 (.A(G5297_1062_gat), .Y(G5303_1417_gat) );
INVXL U_g1218 (.A(G6522_1063_gat), .Y(G6526_1418_gat) );
INVXL U_g1219 (.A(G7327_1064_gat), .Y(G7333_1419_gat) );
INVXL U_g1220 (.A(G6370_1065_gat), .Y(G6374_1420_gat) );
INVXL U_g1221 (.A(G6378_1066_gat), .Y(G6382_1421_gat) );
INVXL U_g1222 (.A(G7330_1067_gat), .Y(G7334_1422_gat) );
INVXL U_g1223 (.A(G7317_1068_gat), .Y(G7323_1423_gat) );
INVXL U_g1224 (.A(G6386_1069_gat), .Y(G6390_1424_gat) );
INVXL U_g1225 (.A(G6426_1070_gat), .Y(G6430_1425_gat) );
INVXL U_g1226 (.A(G7320_1071_gat), .Y(G7324_1426_gat) );
INVXL U_g1227 (.A(G7309_1072_gat), .Y(G7315_1427_gat) );
INVXL U_g1228 (.A(G6394_1073_gat), .Y(G6398_1428_gat) );
INVXL U_g1229 (.A(G5339_1074_gat), .Y(G5345_1429_gat) );
INVXL U_g1230 (.A(G5764_1075_gat), .Y(G5768_1430_gat) );
INVXL U_g1231 (.A(G5412_1076_gat), .Y(G5416_1431_gat) );
INVXL U_g1232 (.A(G5452_1077_gat), .Y(G5456_1432_gat) );
INVXL U_g1233 (.A(G5772_1078_gat), .Y(G5776_1433_gat) );
INVXL U_g1234 (.A(G5342_1079_gat), .Y(G5346_1434_gat) );
INVXL U_g1235 (.A(G5331_1080_gat), .Y(G5337_1435_gat) );
INVXL U_g1236 (.A(G5780_1081_gat), .Y(G5784_1436_gat) );
INVXL U_g1237 (.A(G5420_1082_gat), .Y(G5424_1437_gat) );
INVXL U_g1238 (.A(G5349_1083_gat), .Y(G5355_1438_gat) );
INVXL U_g1239 (.A(G5396_1084_gat), .Y(G5400_1439_gat) );
INVXL U_g1240 (.A(G5748_1085_gat), .Y(G5752_1440_gat) );
INVXL U_g1241 (.A(G5756_1086_gat), .Y(G5760_1441_gat) );
INVXL U_g1242 (.A(G5404_1087_gat), .Y(G5408_1442_gat) );
INVXL U_g1243 (.A(G5352_1088_gat), .Y(G5356_1443_gat) );
INVXL U_g1244 (.A(G5202_1089_gat), .Y(G5206_1444_gat) );
INVXL U_g1245 (.A(G4892_1090_gat), .Y(G4896_1445_gat) );
INVXL U_g1246 (.A(G5266_1091_gat), .Y(G5270_1446_gat) );
INVXL U_g1247 (.A(G5255_1092_gat), .Y(G5261_1447_gat) );
INVXL U_g1248 (.A(G4900_1093_gat), .Y(G4904_1448_gat) );
INVXL U_g1249 (.A(G5210_1094_gat), .Y(G5214_1449_gat) );
INVXL U_g1250 (.A(G5218_1095_gat), .Y(G5222_1450_gat) );
INVXL U_g1251 (.A(G4908_1096_gat), .Y(G4912_1451_gat) );
INVXL U_g1252 (.A(G5258_1097_gat), .Y(G5262_1452_gat) );
INVXL U_g1253 (.A(G5247_1098_gat), .Y(G5253_1453_gat) );
INVXL U_g1254 (.A(G4924_1099_gat), .Y(G4928_1454_gat) );
INVXL U_g1255 (.A(G5226_1100_gat), .Y(G5230_1455_gat) );
INVXL U_g1256 (.A(G5250_1101_gat), .Y(G5254_1456_gat) );
OR2XL U_g1257 (.A(G5278_1103_ngat), .B(G5271_863_ngat), .Y(G5280_1457_gat) );
OR2XL U_g1258 (.A(G5277_1102_ngat), .B(G5274_864_ngat), .Y(G5279_1458_gat) );
INVXL U_g1259 (.A(G5263_1104_gat), .Y(G5269_1459_gat) );
INVXL U_g1260 (.A(G4884_1105_gat), .Y(G4888_1460_gat) );
INVXL U_g1261 (.A(G5194_1106_gat), .Y(G5198_1461_gat) );
AND2XL U_g1262 (.A(G3170_866_gat), .B(G3212_1367_gat), .Y(G3216_1462_gat) );
OR2XL U_g1263 (.A(G6859_431_ngat), .B(G6856_1327_ngat), .Y(G3843_1463_gat) );
OR2XL U_g1264 (.A(G6573_432_ngat), .B(G6570_1329_ngat), .Y(G3281_1464_gat) );
OR2XL U_g1265 (.A(G6581_433_ngat), .B(G6578_1350_ngat), .Y(G3293_1465_gat) );
OR2XL U_g1266 (.A(G6867_434_ngat), .B(G6864_1352_ngat), .Y(G3854_1466_gat) );
OR2XL U_g1267 (.A(G6589_435_ngat), .B(G6586_1378_ngat), .Y(G3312_1467_gat) );
OR2XL U_g1268 (.A(G6875_436_ngat), .B(G6872_1377_ngat), .Y(G3872_1468_gat) );
BUFX20 U_g1269 (.A(G3335_1113_gat), .Y(G6679_1469_gat) );
BUFX20 U_g1270 (.A(G3891_1114_gat), .Y(G6983_1470_gat) );
INVXL U_g1271 (.A(G6925_1115_gat), .Y(G6931_1471_gat) );
OR2XL U_g1272 (.A(G6915_437_ngat), .B(G6912_1374_ngat), .Y(G3987_1472_gat) );
OR2XL U_g1273 (.A(G6597_438_ngat), .B(G6594_1375_ngat), .Y(G3342_1473_gat) );
INVXL U_g1274 (.A(G6671_1116_gat), .Y(G6677_1474_gat) );
OR2XL U_g1275 (.A(G6883_439_ngat), .B(G6880_1361_ngat), .Y(G3897_1475_gat) );
OR2XL U_g1276 (.A(G6605_440_ngat), .B(G6602_1359_ngat), .Y(G3351_1476_gat) );
OR2XL U_g1277 (.A(G6613_441_ngat), .B(G6610_1266_ngat), .Y(G3363_1477_gat) );
OR2XL U_g1278 (.A(G6891_442_ngat), .B(G6888_1267_ngat), .Y(G3909_1478_gat) );
OR2XL U_g1279 (.A(G6899_443_ngat), .B(G6896_1302_ngat), .Y(G3930_1479_gat) );
OR2XL U_g1280 (.A(G6621_444_ngat), .B(G6618_1303_ngat), .Y(G3379_1480_gat) );
OR2XL U_g1281 (.A(G6907_445_ngat), .B(G6904_1296_ngat), .Y(G3955_1481_gat) );
OR2XL U_g1282 (.A(G6629_446_ngat), .B(G6626_1297_ngat), .Y(G3397_1482_gat) );
BUFX20 U_g1283 (.A(G3979_1126_gat), .Y(G7129_1483_gat) );
OR2XL U_g1284 (.A(G6637_447_ngat), .B(G6634_1275_ngat), .Y(G3415_1484_gat) );
INVXL U_g1285 (.A(G7041_1127_gat), .Y(G7047_1485_gat) );
OR2XL U_g1286 (.A(G6923_448_ngat), .B(G6920_1276_ngat), .Y(G3995_1486_gat) );
OR2XL U_g1287 (.A(G5991_449_ngat), .B(G5988_1290_ngat), .Y(G2587_1487_gat) );
OR2XL U_g1288 (.A(G5871_450_ngat), .B(G5868_1291_ngat), .Y(G2341_1488_gat) );
OR2XL U_g1289 (.A(G5879_451_ngat), .B(G5876_1259_ngat), .Y(G2352_1489_gat) );
OR2XL U_g1290 (.A(G5999_452_ngat), .B(G5996_1260_ngat), .Y(G2598_1490_gat) );
OR2XL U_g1291 (.A(G6007_453_ngat), .B(G6004_1254_ngat), .Y(G2616_1491_gat) );
OR2XL U_g1292 (.A(G5887_454_ngat), .B(G5884_1255_ngat), .Y(G2370_1492_gat) );
BUFX20 U_g1293 (.A(G2391_1134_gat), .Y(G5977_1493_gat) );
BUFX20 U_g1294 (.A(G2635_1135_gat), .Y(G6115_1494_gat) );
INVXL U_g1295 (.A(G6057_1136_gat), .Y(G6063_1495_gat) );
OR2XL U_g1296 (.A(G6047_455_ngat), .B(G6044_1251_ngat), .Y(G2732_1496_gat) );
OR2XL U_g1297 (.A(G5895_456_ngat), .B(G5892_1250_ngat), .Y(G2398_1497_gat) );
INVXL U_g1298 (.A(G5969_1137_gat), .Y(G5975_1498_gat) );
OR2XL U_g1299 (.A(G5903_457_ngat), .B(G5900_1288_ngat), .Y(G2407_1499_gat) );
OR2XL U_g1300 (.A(G6015_458_ngat), .B(G6012_1287_ngat), .Y(G2641_1500_gat) );
OR2XL U_g1301 (.A(G6023_459_ngat), .B(G6020_1395_ngat), .Y(G2653_1501_gat) );
OR2XL U_g1302 (.A(G5911_460_ngat), .B(G5908_1394_ngat), .Y(G2418_1502_gat) );
OR2XL U_g1303 (.A(G5919_461_ngat), .B(G5916_1390_ngat), .Y(G2434_1503_gat) );
OR2XL U_g1304 (.A(G6031_462_ngat), .B(G6028_1389_ngat), .Y(G2674_1504_gat) );
OR2XL U_g1305 (.A(G6039_463_ngat), .B(G6036_1383_ngat), .Y(G2699_1505_gat) );
OR2XL U_g1306 (.A(G5927_464_ngat), .B(G5924_1382_ngat), .Y(G2452_1506_gat) );
OR2XL U_g1307 (.A(G7504_1150_ngat), .B(G7497_868_ngat), .Y(G7506_1507_gat) );
OR2XL U_g1308 (.A(G6374_1420_ngat), .B(G6367_869_ngat), .Y(G2955_1508_gat) );
OR2XL U_g1309 (.A(G5400_1439_ngat), .B(G5393_352_ngat), .Y(G1545_1509_gat) );
OR2XL U_g1310 (.A(G5752_1440_ngat), .B(G5745_353_ngat), .Y(G1794_1510_gat) );
OR2XL U_g1311 (.A(G7503_1146_ngat), .B(G7500_873_ngat), .Y(G7505_1511_gat) );
OR2XL U_g1312 (.A(G6382_1421_ngat), .B(G6375_874_ngat), .Y(G2964_1512_gat) );
OR2XL U_g1313 (.A(G5760_1441_ngat), .B(G5753_354_ngat), .Y(G1804_1513_gat) );
OR2XL U_g1314 (.A(G5408_1442_ngat), .B(G5401_355_ngat), .Y(G1555_1514_gat) );
OR2XL U_g1315 (.A(G6390_1424_ngat), .B(G6383_880_ngat), .Y(G2972_1515_gat) );
OR2XL U_g1316 (.A(G7494_1164_ngat), .B(G7487_881_ngat), .Y(G7496_1516_gat) );
OR2XL U_g1317 (.A(G5416_1431_ngat), .B(G5409_356_ngat), .Y(G1572_1517_gat) );
OR2XL U_g1318 (.A(G5768_1430_ngat), .B(G5761_357_ngat), .Y(G1821_1518_gat) );
INVXL U_g1319 (.A(G5523_1158_gat), .Y(G5529_1519_gat) );
INVXL U_g1320 (.A(G5857_1159_gat), .Y(G5863_1520_gat) );
OR2XL U_g1321 (.A(G5776_1433_ngat), .B(G5769_358_ngat), .Y(G1849_1521_gat) );
OR2XL U_g1322 (.A(G5456_1432_ngat), .B(G5449_359_ngat), .Y(G1686_1522_gat) );
OR2XL U_g1323 (.A(G7493_1155_ngat), .B(G7490_887_ngat), .Y(G7495_1523_gat) );
OR2XL U_g1324 (.A(G6430_1425_ngat), .B(G6423_888_ngat), .Y(G3017_1524_gat) );
OR2XL U_g1325 (.A(G7486_1173_ngat), .B(G7479_890_ngat), .Y(G4548_1525_gat) );
OR2XL U_g1326 (.A(G6398_1428_ngat), .B(G6391_891_ngat), .Y(G2981_1526_gat) );
OR2XL U_g1327 (.A(G5424_1437_ngat), .B(G5417_360_ngat), .Y(G1597_1527_gat) );
OR2XL U_g1328 (.A(G5784_1436_ngat), .B(G5777_361_ngat), .Y(G1858_1528_gat) );
OR2XL U_g1329 (.A(G5792_1243_ngat), .B(G5785_362_ngat), .Y(G1868_1529_gat) );
OR2XL U_g1330 (.A(G5432_1242_ngat), .B(G5425_363_ngat), .Y(G1608_1530_gat) );
OR2XL U_g1331 (.A(G6406_1230_ngat), .B(G6399_897_ngat), .Y(G2991_1531_gat) );
OR2XL U_g1332 (.A(G7485_1166_ngat), .B(G7482_898_ngat), .Y(G4547_1532_gat) );
OR2XL U_g1333 (.A(G7478_1181_ngat), .B(G7471_902_ngat), .Y(G4539_1533_gat) );
OR2XL U_g1334 (.A(G6414_1229_ngat), .B(G6407_903_ngat), .Y(G3000_1534_gat) );
OR2XL U_g1335 (.A(G5440_1240_ngat), .B(G5433_364_ngat), .Y(G1629_1535_gat) );
OR2XL U_g1336 (.A(G5800_1239_ngat), .B(G5793_365_ngat), .Y(G1884_1536_gat) );
OR2XL U_g1337 (.A(G5808_1237_ngat), .B(G5801_366_ngat), .Y(G1902_1537_gat) );
OR2XL U_g1338 (.A(G5448_1236_ngat), .B(G5441_367_ngat), .Y(G1654_1538_gat) );
OR2XL U_g1339 (.A(G6422_1226_ngat), .B(G6415_907_ngat), .Y(G3008_1539_gat) );
OR2XL U_g1340 (.A(G7477_1174_ngat), .B(G7474_908_ngat), .Y(G4538_1540_gat) );
INVXL U_g1341 (.A(G5669_1182_gat), .Y(G5675_1541_gat) );
OR2XL U_g1342 (.A(G5464_1246_ngat), .B(G5457_368_ngat), .Y(G1694_1542_gat) );
OR2XL U_g1343 (.A(G6438_1233_ngat), .B(G6431_914_ngat), .Y(G3020_1543_gat) );
OR2XL U_g1344 (.A(G5816_1245_ngat), .B(G5809_369_ngat), .Y(G1920_1544_gat) );
OR2XL U_g1345 (.A(G7469_1186_ngat), .B(G7466_771_ngat), .Y(G4529_1545_gat) );
OR2XL U_g1346 (.A(G6720_1189_ngat), .B(G6719_1202_ngat), .Y(G6832_1546_gat) );
OR2XL U_g1347 (.A(G953_1197_gat), .B(G917_1190_gat), .Y(G4932_1547_gat) );
INVXL U_g1348 (.A(G917_1190_gat), .Y(G4973_1548_gat) );
INVXL U_g1349 (.A(G4983_1191_gat), .Y(G4987_1549_gat) );
INVXL U_g1350 (.A(G908_1192_gat), .Y(G912_1550_gat) );
OR3XL U_g1351 (.A(G914_1200_gat), .B(G913_1027_gat), .C(G777_370_gat), .Y(G4942_1551_gat) );
INVXL U_g1352 (.A(G1117_1193_gat), .Y(G1121_1552_gat) );
INVXL U_g1353 (.A(G1108_1196_gat), .Y(G1112_1553_gat) );
INVXL U_g1354 (.A(G902_1199_gat), .Y(G906_1554_gat) );
INVXL U_g1355 (.A(G4993_1203_gat), .Y(G4997_1555_gat) );
INVXL U_g1356 (.A(G4952_1204_gat), .Y(G4956_1556_gat) );
OR2XL U_g1357 (.A(G6710_1213_ngat), .B(G6703_927_ngat), .Y(G3521_1557_gat) );
OR2XL U_g1358 (.A(G6526_1418_ngat), .B(G6519_928_ngat), .Y(G3175_1558_gat) );
OR2XL U_g1359 (.A(G4888_1460_ngat), .B(G4881_375_ngat), .Y(G791_1559_gat) );
OR2XL U_g1360 (.A(G5198_1461_ngat), .B(G5191_376_ngat), .Y(G1025_1560_gat) );
OR2XL U_g1361 (.A(G5206_1444_ngat), .B(G5199_377_ngat), .Y(G1037_1561_gat) );
OR2XL U_g1362 (.A(G4896_1445_ngat), .B(G4889_378_ngat), .Y(G804_1562_gat) );
OR2XL U_g1363 (.A(G6534_1408_ngat), .B(G6527_932_ngat), .Y(G3185_1563_gat) );
OR2XL U_g1364 (.A(G6709_1206_ngat), .B(G6706_933_ngat), .Y(G3520_1564_gat) );
OR2XL U_g1365 (.A(G5222_1450_ngat), .B(G5215_379_ngat), .Y(G1073_1565_gat) );
OR2XL U_g1366 (.A(G6550_1412_ngat), .B(G6543_937_ngat), .Y(G3202_1566_gat) );
OR2XL U_g1367 (.A(G6701_1281_ngat), .B(G6698_938_ngat), .Y(G3511_1567_gat) );
OR2XL U_g1368 (.A(G4912_1451_ngat), .B(G4905_380_ngat), .Y(G852_1568_gat) );
INVXL U_g1369 (.A(G5099_1218_gat), .Y(G5105_1569_gat) );
OR2XL U_g1370 (.A(G4928_1454_ngat), .B(G4921_381_ngat), .Y(G894_1570_gat) );
OR2XL U_g1371 (.A(G6566_1414_ngat), .B(G6559_944_ngat), .Y(G3214_1571_gat) );
OR2XL U_g1372 (.A(G5230_1455_ngat), .B(G5223_382_ngat), .Y(G1092_1572_gat) );
OR2XL U_g1373 (.A(G6693_1222_ngat), .B(G6690_780_ngat), .Y(G3502_1573_gat) );
OR2XL U_g1374 (.A(G7299_1232_ngat), .B(G7296_811_ngat), .Y(G4224_1574_gat) );
OR2XL U_g1375 (.A(G6421_1180_ngat), .B(G6418_947_ngat), .Y(G3007_1575_gat) );
OR2XL U_g1376 (.A(G7307_1228_ngat), .B(G7304_948_ngat), .Y(G4233_1576_gat) );
OR2XL U_g1377 (.A(G7308_1227_ngat), .B(G7301_949_ngat), .Y(G4234_1577_gat) );
OR2XL U_g1378 (.A(G6413_1175_ngat), .B(G6410_950_ngat), .Y(G2999_1578_gat) );
OR2XL U_g1379 (.A(G6405_1172_ngat), .B(G6402_951_ngat), .Y(G2990_1579_gat) );
OR2XL U_g1380 (.A(G7315_1427_ngat), .B(G7312_952_ngat), .Y(G4242_1580_gat) );
OR2XL U_g1381 (.A(G6437_1187_ngat), .B(G6434_954_ngat), .Y(G3019_1581_gat) );
OR2XL U_g1382 (.A(G5321_1244_ngat), .B(G5318_816_ngat), .Y(G1261_1582_gat) );
OR2XL U_g1383 (.A(G5329_1238_ngat), .B(G5326_956_ngat), .Y(G1270_1583_gat) );
OR2XL U_g1384 (.A(G5330_1235_ngat), .B(G5323_959_ngat), .Y(G1271_1584_gat) );
OR2XL U_g1385 (.A(G5337_1435_ngat), .B(G5334_962_ngat), .Y(G1279_1585_gat) );
INVXL U_g1386 (.A(G7276_1247_gat), .Y(G7280_1586_gat) );
INVXL U_g1387 (.A(G7420_1249_gat), .Y(G7424_1587_gat) );
INVXL U_g1388 (.A(G5892_1250_gat), .Y(G5896_1588_gat) );
INVXL U_g1389 (.A(G6044_1251_gat), .Y(G6048_1589_gat) );
INVXL U_g1390 (.A(G6792_1252_gat), .Y(G6796_1590_gat) );
INVXL U_g1391 (.A(G6789_1253_gat), .Y(G6795_1591_gat) );
INVXL U_g1392 (.A(G6004_1254_gat), .Y(G6008_1592_gat) );
INVXL U_g1393 (.A(G5884_1255_gat), .Y(G5888_1593_gat) );
INVXL U_g1394 (.A(G7380_1257_gat), .Y(G7384_1594_gat) );
INVXL U_g1395 (.A(G7273_1258_gat), .Y(G7279_1595_gat) );
INVXL U_g1396 (.A(G5876_1259_gat), .Y(G5880_1596_gat) );
INVXL U_g1397 (.A(G5996_1260_gat), .Y(G6000_1597_gat) );
INVXL U_g1398 (.A(G6802_1261_gat), .Y(G6806_1598_gat) );
INVXL U_g1399 (.A(G7372_1263_gat), .Y(G7376_1599_gat) );
INVXL U_g1400 (.A(G7286_1264_gat), .Y(G7290_1600_gat) );
INVXL U_g1401 (.A(G6740_1265_gat), .Y(G6744_1601_gat) );
INVXL U_g1402 (.A(G6610_1266_gat), .Y(G6614_1602_gat) );
INVXL U_g1403 (.A(G6888_1267_gat), .Y(G6892_1603_gat) );
INVXL U_g1404 (.A(G6474_1269_gat), .Y(G6478_1604_gat) );
OR2XL U_g1405 (.A(G7227_1358_ngat), .B(G7224_1270_ngat), .Y(G4196_1605_gat) );
INVXL U_g1406 (.A(G7224_1270_gat), .Y(G7228_1606_gat) );
INVXL U_g1407 (.A(G6506_1272_gat), .Y(G6510_1607_gat) );
OR2XL U_g1408 (.A(G7212_1277_ngat), .B(G7205_1273_ngat), .Y(G4179_1608_gat) );
INVXL U_g1409 (.A(G7205_1273_gat), .Y(G7211_1609_gat) );
OR2XL U_g1410 (.A(G6728_1278_ngat), .B(G6721_1274_ngat), .Y(G3526_1610_gat) );
INVXL U_g1411 (.A(G6721_1274_gat), .Y(G6727_1611_gat) );
INVXL U_g1412 (.A(G6634_1275_gat), .Y(G6638_1612_gat) );
INVXL U_g1413 (.A(G6920_1276_gat), .Y(G6924_1613_gat) );
OR2XL U_g1414 (.A(G4904_1448_ngat), .B(G4897_548_ngat), .Y(G826_1614_gat) );
OR2XL U_g1415 (.A(G5214_1449_ngat), .B(G5207_549_ngat), .Y(G1054_1615_gat) );
OR2XL U_g1416 (.A(G6702_1216_ngat), .B(G6695_983_ngat), .Y(G3512_1616_gat) );
OR2XL U_g1417 (.A(G6542_1410_ngat), .B(G6535_984_ngat), .Y(G3194_1617_gat) );
INVXL U_g1418 (.A(G7388_1283_gat), .Y(G7392_1618_gat) );
OR2XL U_g1419 (.A(G7272_1399_ngat), .B(G7265_1285_ngat), .Y(G4220_1619_gat) );
INVXL U_g1420 (.A(G7265_1285_gat), .Y(G7271_1620_gat) );
INVXL U_g1421 (.A(G6781_1286_gat), .Y(G6787_1621_gat) );
INVXL U_g1422 (.A(G6012_1287_gat), .Y(G6016_1622_gat) );
INVXL U_g1423 (.A(G5900_1288_gat), .Y(G5904_1623_gat) );
INVXL U_g1424 (.A(G6799_1289_gat), .Y(G6805_1624_gat) );
INVXL U_g1425 (.A(G5988_1290_gat), .Y(G5992_1625_gat) );
INVXL U_g1426 (.A(G5868_1291_gat), .Y(G5872_1626_gat) );
INVXL U_g1427 (.A(G7364_1292_gat), .Y(G7368_1627_gat) );
INVXL U_g1428 (.A(G7283_1294_gat), .Y(G7289_1628_gat) );
INVXL U_g1429 (.A(G6732_1295_gat), .Y(G6736_1629_gat) );
INVXL U_g1430 (.A(G6904_1296_gat), .Y(G6908_1630_gat) );
INVXL U_g1431 (.A(G6626_1297_gat), .Y(G6630_1631_gat) );
INVXL U_g1432 (.A(G6490_1299_gat), .Y(G6494_1632_gat) );
INVXL U_g1433 (.A(G7216_1300_gat), .Y(G7220_1633_gat) );
INVXL U_g1434 (.A(G6729_1301_gat), .Y(G6735_1634_gat) );
INVXL U_g1435 (.A(G6896_1302_gat), .Y(G6900_1635_gat) );
INVXL U_g1436 (.A(G6618_1303_gat), .Y(G6622_1636_gat) );
INVXL U_g1437 (.A(G6482_1304_gat), .Y(G6486_1637_gat) );
INVXL U_g1438 (.A(G7213_1306_gat), .Y(G7219_1638_gat) );
INVXL U_g1439 (.A(G6471_1307_gat), .Y(G6477_1639_gat) );
INVXL U_g1440 (.A(G7570_1308_gat), .Y(G7574_1640_gat) );
OR2XL U_g1441 (.A(G6470_1357_ngat), .B(G6463_1309_ngat), .Y(G3081_1641_gat) );
INVXL U_g1442 (.A(G6463_1309_gat), .Y(G6469_1642_gat) );
INVXL U_g1443 (.A(G7567_1310_gat), .Y(G7573_1643_gat) );
OR2XL U_g1444 (.A(G6502_1371_ngat), .B(G6495_1311_ngat), .Y(G3118_1644_gat) );
INVXL U_g1445 (.A(G6495_1311_gat), .Y(G6501_1645_gat) );
INVXL U_g1446 (.A(G7578_1312_gat), .Y(G7582_1646_gat) );
INVXL U_g1447 (.A(G6487_1313_gat), .Y(G6493_1647_gat) );
INVXL U_g1448 (.A(G7562_1314_gat), .Y(G7566_1648_gat) );
INVXL U_g1449 (.A(G6503_1315_gat), .Y(G6509_1649_gat) );
OR2XL U_g1450 (.A(G7558_1341_ngat), .B(G7551_1316_ngat), .Y(G4576_1650_gat) );
INVXL U_g1451 (.A(G7551_1316_gat), .Y(G7557_1651_gat) );
INVXL U_g1452 (.A(G7515_1317_gat), .Y(G7521_1652_gat) );
OR2XL U_g1453 (.A(G7408_1391_ngat), .B(G7401_1318_ngat), .Y(G4335_1653_gat) );
INVXL U_g1454 (.A(G7401_1318_gat), .Y(G7407_1654_gat) );
OR2XL U_g1455 (.A(G7400_1398_ngat), .B(G7393_1319_ngat), .Y(G4326_1655_gat) );
INVXL U_g1456 (.A(G7393_1319_gat), .Y(G7399_1656_gat) );
INVXL U_g1457 (.A(G7526_1320_gat), .Y(G7530_1657_gat) );
OR2XL U_g1458 (.A(G7416_1386_ngat), .B(G7409_1321_ngat), .Y(G4343_1658_gat) );
INVXL U_g1459 (.A(G7409_1321_gat), .Y(G7415_1659_gat) );
INVXL U_g1460 (.A(G7518_1322_gat), .Y(G7522_1660_gat) );
INVXL U_g1461 (.A(G7523_1323_gat), .Y(G7529_1661_gat) );
INVXL U_g1462 (.A(G7385_1324_gat), .Y(G7391_1662_gat) );
OR2XL U_g1463 (.A(G7514_1326_ngat), .B(G7507_1002_ngat), .Y(G4553_1663_gat) );
OR2XL U_g1464 (.A(G7513_1325_ngat), .B(G7510_1003_ngat), .Y(G4552_1664_gat) );
INVXL U_g1465 (.A(G6856_1327_gat), .Y(G6860_1665_gat) );
INVXL U_g1466 (.A(G6755_1328_gat), .Y(G6761_1666_gat) );
INVXL U_g1467 (.A(G6570_1329_gat), .Y(G6574_1667_gat) );
OR2XL U_g1468 (.A(G7246_1355_ngat), .B(G7239_1005_ngat), .Y(G7248_1668_gat) );
OR2XL U_g1469 (.A(G6446_1332_ngat), .B(G6439_1333_ngat), .Y(G3051_1669_gat) );
INVXL U_g1470 (.A(G6439_1333_gat), .Y(G6445_1670_gat) );
INVXL U_g1471 (.A(G7585_1334_gat), .Y(G7591_1671_gat) );
OR2XL U_g1472 (.A(G6454_1354_ngat), .B(G6447_1335_ngat), .Y(G3061_1672_gat) );
INVXL U_g1473 (.A(G6447_1335_gat), .Y(G6453_1673_gat) );
INVXL U_g1474 (.A(G7588_1336_gat), .Y(G7592_1674_gat) );
OR2XL U_g1475 (.A(G6462_1380_ngat), .B(G6455_1337_ngat), .Y(G3070_1675_gat) );
INVXL U_g1476 (.A(G6455_1337_gat), .Y(G6461_1676_gat) );
INVXL U_g1477 (.A(G7575_1338_gat), .Y(G7581_1677_gat) );
INVXL U_g1478 (.A(G6479_1339_gat), .Y(G6485_1678_gat) );
INVXL U_g1479 (.A(G7559_1340_gat), .Y(G7565_1679_gat) );
INVXL U_g1480 (.A(G7541_1342_gat), .Y(G7547_1680_gat) );
INVXL U_g1481 (.A(G7361_1343_gat), .Y(G7367_1681_gat) );
INVXL U_g1482 (.A(G7369_1344_gat), .Y(G7375_1682_gat) );
INVXL U_g1483 (.A(G7544_1345_gat), .Y(G7548_1683_gat) );
INVXL U_g1484 (.A(G7531_1346_gat), .Y(G7537_1684_gat) );
INVXL U_g1485 (.A(G7377_1347_gat), .Y(G7383_1685_gat) );
INVXL U_g1486 (.A(G7534_1348_gat), .Y(G7538_1686_gat) );
INVXL U_g1487 (.A(G7417_1349_gat), .Y(G7423_1687_gat) );
INVXL U_g1488 (.A(G6578_1350_gat), .Y(G6582_1688_gat) );
INVXL U_g1489 (.A(G6758_1351_gat), .Y(G6762_1689_gat) );
INVXL U_g1490 (.A(G6864_1352_gat), .Y(G6868_1690_gat) );
OR2XL U_g1491 (.A(G7245_1331_ngat), .B(G7242_1018_ngat), .Y(G7247_1691_gat) );
INVXL U_g1492 (.A(G6602_1359_gat), .Y(G6606_1692_gat) );
INVXL U_g1493 (.A(G6737_1360_gat), .Y(G6743_1693_gat) );
INVXL U_g1494 (.A(G6880_1361_gat), .Y(G6884_1694_gat) );
OR2XL U_g1495 (.A(G7255_1364_ngat), .B(G7252_825_ngat), .Y(G4201_1695_gat) );
OR2XL U_g1496 (.A(G6772_1363_ngat), .B(G6765_1365_ngat), .Y(G3549_1696_gat) );
INVXL U_g1497 (.A(G6765_1365_gat), .Y(G6771_1697_gat) );
OR2XL U_g1498 (.A(G3222_1366_gat), .B(G3221_557_gat), .Y(G3223_1698_gat) );
OR2XL U_g1499 (.A(G5246_1194_ngat), .B(G5239_719_ngat), .Y(G1157_1699_gat) );
OR2XL U_g1500 (.A(G5238_1195_ngat), .B(G5231_561_ngat), .Y(G1153_1700_gat) );
OR2XL U_g1501 (.A(G7235_1381_ngat), .B(G7232_1033_ngat), .Y(G7237_1701_gat) );
INVXL U_g1502 (.A(G6748_1373_gat), .Y(G6752_1702_gat) );
INVXL U_g1503 (.A(G6912_1374_gat), .Y(G6916_1703_gat) );
INVXL U_g1504 (.A(G6594_1375_gat), .Y(G6598_1704_gat) );
INVXL U_g1505 (.A(G6745_1376_gat), .Y(G6751_1705_gat) );
INVXL U_g1506 (.A(G6872_1377_gat), .Y(G6876_1706_gat) );
INVXL U_g1507 (.A(G6586_1378_gat), .Y(G6590_1707_gat) );
OR2XL U_g1508 (.A(G7236_1372_ngat), .B(G7229_1037_ngat), .Y(G7238_1708_gat) );
INVXL U_g1509 (.A(G5924_1382_gat), .Y(G5928_1709_gat) );
INVXL U_g1510 (.A(G6036_1383_gat), .Y(G6040_1710_gat) );
INVXL U_g1511 (.A(G6776_1384_gat), .Y(G6780_1711_gat) );
OR2XL U_g1512 (.A(G7263_1393_ngat), .B(G7260_1040_ngat), .Y(G4210_1712_gat) );
INVXL U_g1513 (.A(G6773_1388_gat), .Y(G6779_1713_gat) );
INVXL U_g1514 (.A(G6028_1389_gat), .Y(G6032_1714_gat) );
INVXL U_g1515 (.A(G5916_1390_gat), .Y(G5920_1715_gat) );
OR2XL U_g1516 (.A(G7264_1387_ngat), .B(G7257_1043_ngat), .Y(G4211_1716_gat) );
INVXL U_g1517 (.A(G5908_1394_gat), .Y(G5912_1717_gat) );
INVXL U_g1518 (.A(G6020_1395_gat), .Y(G6024_1718_gat) );
INVXL U_g1519 (.A(G6784_1396_gat), .Y(G6788_1719_gat) );
OR2XL U_g1520 (.A(G7431_1401_ngat), .B(G7428_1404_ngat), .Y(G4353_1720_gat) );
AND2XL U_g1521 (.A(G4389_1405_gat), .B(G3682_839_gat), .Y(G2481_1721_gat) );
AND2XL U_g1522 (.A(G4389_1405_gat), .B(G3682_839_gat), .Y(G2724_1722_gat) );
AND2XL U_g1523 (.A(G4389_1405_ngat), .B(G3682_839_ngat), .Y(G6173_1723_gat) );
INVXL U_g1524 (.A(G7428_1404_gat), .Y(G7432_1724_gat) );
BUFX20 U_g1525 (.A(G4389_1405_gat), .Y(G6052_1725_gat) );
BUFX20 U_g1526 (.A(G4389_1405_gat), .Y(G5932_1726_gat) );
OR2XL U_g1527 (.A(G5287_1413_ngat), .B(G5284_1051_ngat), .Y(G1238_1727_gat) );
OR2XL U_g1528 (.A(G5303_1417_ngat), .B(G5300_1052_ngat), .Y(G1256_1728_gat) );
OR2XL U_g1529 (.A(G6533_1212_ngat), .B(G6530_1053_ngat), .Y(G3184_1729_gat) );
OR2XL U_g1530 (.A(G5296_1411_ngat), .B(G5289_1054_ngat), .Y(G1248_1730_gat) );
OR2XL U_g1531 (.A(G6541_1282_ngat), .B(G6538_1055_ngat), .Y(G3193_1731_gat) );
OR2XL U_g1532 (.A(G5295_1409_ngat), .B(G5292_1056_ngat), .Y(G1247_1732_gat) );
OR2XL U_g1533 (.A(G6549_1215_ngat), .B(G6546_1057_ngat), .Y(G3201_1733_gat) );
OR2XL U_g1534 (.A(G5288_1406_ngat), .B(G5281_1058_ngat), .Y(G1239_1734_gat) );
OR2XL U_g1535 (.A(G6565_1223_ngat), .B(G6562_1059_ngat), .Y(G3213_1735_gat) );
OR2XL U_g1536 (.A(G5314_1415_ngat), .B(G5313_1416_ngat), .Y(G5380_1736_gat) );
OR2XL U_g1537 (.A(G5304_1407_ngat), .B(G5297_1062_ngat), .Y(G1257_1737_gat) );
OR2XL U_g1538 (.A(G6525_1207_ngat), .B(G6522_1063_ngat), .Y(G3174_1738_gat) );
OR2XL U_g1539 (.A(G7334_1422_ngat), .B(G7327_1064_ngat), .Y(G7336_1739_gat) );
OR2XL U_g1540 (.A(G6373_1147_ngat), .B(G6370_1065_ngat), .Y(G2954_1740_gat) );
OR2XL U_g1541 (.A(G6381_1151_ngat), .B(G6378_1066_ngat), .Y(G2963_1741_gat) );
OR2XL U_g1542 (.A(G7333_1419_ngat), .B(G7330_1067_ngat), .Y(G7335_1742_gat) );
OR2XL U_g1543 (.A(G7324_1426_ngat), .B(G7317_1068_ngat), .Y(G7326_1743_gat) );
OR2XL U_g1544 (.A(G6389_1154_ngat), .B(G6386_1069_ngat), .Y(G2971_1744_gat) );
OR2XL U_g1545 (.A(G6429_1165_ngat), .B(G6426_1070_ngat), .Y(G3016_1745_gat) );
OR2XL U_g1546 (.A(G7323_1423_ngat), .B(G7320_1071_ngat), .Y(G7325_1746_gat) );
OR2XL U_g1547 (.A(G7316_1231_ngat), .B(G7309_1072_ngat), .Y(G4243_1747_gat) );
OR2XL U_g1548 (.A(G6397_1167_ngat), .B(G6394_1073_ngat), .Y(G2980_1748_gat) );
OR2XL U_g1549 (.A(G5346_1434_ngat), .B(G5339_1074_ngat), .Y(G5348_1749_gat) );
OR2XL U_g1550 (.A(G5345_1429_ngat), .B(G5342_1079_ngat), .Y(G5347_1750_gat) );
OR2XL U_g1551 (.A(G5338_1241_ngat), .B(G5331_1080_ngat), .Y(G1280_1751_gat) );
OR2XL U_g1552 (.A(G5356_1443_ngat), .B(G5349_1083_ngat), .Y(G5358_1752_gat) );
OR2XL U_g1553 (.A(G5355_1438_ngat), .B(G5352_1088_ngat), .Y(G5357_1753_gat) );
OR2XL U_g1554 (.A(G5269_1459_ngat), .B(G5266_1091_ngat), .Y(G1233_1754_gat) );
OR2XL U_g1555 (.A(G5262_1452_ngat), .B(G5255_1092_ngat), .Y(G1225_1755_gat) );
OR2XL U_g1556 (.A(G5261_1447_ngat), .B(G5258_1097_ngat), .Y(G1224_1756_gat) );
OR2XL U_g1557 (.A(G5254_1456_ngat), .B(G5247_1098_ngat), .Y(G1216_1757_gat) );
OR2XL U_g1558 (.A(G5253_1453_ngat), .B(G5250_1101_ngat), .Y(G1215_1758_gat) );
OR2XL U_g1559 (.A(G5280_1457_ngat), .B(G5279_1458_ngat), .Y(G5372_1759_gat) );
OR2XL U_g1560 (.A(G5270_1446_ngat), .B(G5263_1104_ngat), .Y(G1234_1760_gat) );
INVXL U_g1561 (.A(G3216_1462_gat), .Y(G3220_1761_gat) );
OR2XL U_g1562 (.A(G6860_1665_ngat), .B(G6853_318_ngat), .Y(G3844_1762_gat) );
OR2XL U_g1563 (.A(G6574_1667_ngat), .B(G6567_319_ngat), .Y(G3282_1763_gat) );
OR2XL U_g1564 (.A(G6582_1688_ngat), .B(G6575_320_ngat), .Y(G3294_1764_gat) );
OR2XL U_g1565 (.A(G6868_1690_ngat), .B(G6861_321_ngat), .Y(G3855_1765_gat) );
OR2XL U_g1566 (.A(G6590_1707_ngat), .B(G6583_322_ngat), .Y(G3313_1766_gat) );
OR2XL U_g1567 (.A(G6876_1706_ngat), .B(G6869_323_ngat), .Y(G3873_1767_gat) );
INVXL U_g1568 (.A(G6679_1469_gat), .Y(G6685_1768_gat) );
INVXL U_g1569 (.A(G6983_1470_gat), .Y(G6989_1769_gat) );
OR2XL U_g1570 (.A(G6916_1703_ngat), .B(G6909_324_ngat), .Y(G3988_1770_gat) );
OR2XL U_g1571 (.A(G6598_1704_ngat), .B(G6591_325_ngat), .Y(G3343_1771_gat) );
OR2XL U_g1572 (.A(G6884_1694_ngat), .B(G6877_326_ngat), .Y(G3898_1772_gat) );
OR2XL U_g1573 (.A(G6606_1692_ngat), .B(G6599_327_ngat), .Y(G3352_1773_gat) );
OR2XL U_g1574 (.A(G6614_1602_ngat), .B(G6607_328_ngat), .Y(G3364_1774_gat) );
OR2XL U_g1575 (.A(G6892_1603_ngat), .B(G6885_329_ngat), .Y(G3910_1775_gat) );
OR2XL U_g1576 (.A(G6900_1635_ngat), .B(G6893_330_ngat), .Y(G3931_1776_gat) );
OR2XL U_g1577 (.A(G6622_1636_ngat), .B(G6615_331_ngat), .Y(G3380_1777_gat) );
OR2XL U_g1578 (.A(G6908_1630_ngat), .B(G6901_332_ngat), .Y(G3956_1778_gat) );
OR2XL U_g1579 (.A(G6630_1631_ngat), .B(G6623_333_ngat), .Y(G3398_1779_gat) );
INVXL U_g1580 (.A(G7129_1483_gat), .Y(G7135_1780_gat) );
OR2XL U_g1581 (.A(G6638_1612_ngat), .B(G6631_334_ngat), .Y(G3416_1781_gat) );
OR2XL U_g1582 (.A(G6924_1613_ngat), .B(G6917_335_ngat), .Y(G3996_1782_gat) );
OR2XL U_g1583 (.A(G5992_1625_ngat), .B(G5985_336_ngat), .Y(G2588_1783_gat) );
OR2XL U_g1584 (.A(G5872_1626_ngat), .B(G5865_337_ngat), .Y(G2342_1784_gat) );
OR2XL U_g1585 (.A(G5880_1596_ngat), .B(G5873_338_ngat), .Y(G2353_1785_gat) );
OR2XL U_g1586 (.A(G6000_1597_ngat), .B(G5993_339_ngat), .Y(G2599_1786_gat) );
OR2XL U_g1587 (.A(G6008_1592_ngat), .B(G6001_340_ngat), .Y(G2617_1787_gat) );
OR2XL U_g1588 (.A(G5888_1593_ngat), .B(G5881_341_ngat), .Y(G2371_1788_gat) );
INVXL U_g1589 (.A(G5977_1493_gat), .Y(G5983_1789_gat) );
INVXL U_g1590 (.A(G6115_1494_gat), .Y(G6121_1790_gat) );
OR2XL U_g1591 (.A(G6048_1589_ngat), .B(G6041_342_ngat), .Y(G2733_1791_gat) );
OR2XL U_g1592 (.A(G5896_1588_ngat), .B(G5889_343_ngat), .Y(G2399_1792_gat) );
OR2XL U_g1593 (.A(G5904_1623_ngat), .B(G5897_344_ngat), .Y(G2408_1793_gat) );
OR2XL U_g1594 (.A(G6016_1622_ngat), .B(G6009_345_ngat), .Y(G2642_1794_gat) );
OR2XL U_g1595 (.A(G6024_1718_ngat), .B(G6017_346_ngat), .Y(G2654_1795_gat) );
OR2XL U_g1596 (.A(G5912_1717_ngat), .B(G5905_347_ngat), .Y(G2419_1796_gat) );
OR2XL U_g1597 (.A(G5920_1715_ngat), .B(G5913_348_ngat), .Y(G2435_1797_gat) );
OR2XL U_g1598 (.A(G6032_1714_ngat), .B(G6025_349_ngat), .Y(G2675_1798_gat) );
OR2XL U_g1599 (.A(G6040_1710_ngat), .B(G6033_350_ngat), .Y(G2700_1799_gat) );
OR2XL U_g1600 (.A(G5928_1709_ngat), .B(G5921_351_ngat), .Y(G2453_1800_gat) );
OR2XL U_g1601 (.A(G7506_1507_ngat), .B(G7505_1511_ngat), .Y(G7595_1801_gat) );
OR2XL U_g1602 (.A(G2955_1508_ngat), .B(G2954_1740_ngat), .Y(G2956_1802_gat) );
OR2XL U_g1603 (.A(G1545_1509_ngat), .B(G1544_1148_ngat), .Y(G1546_1803_gat) );
OR2XL U_g1604 (.A(G1794_1510_ngat), .B(G1793_1149_ngat), .Y(G1795_1804_gat) );
OR2XL U_g1605 (.A(G2964_1512_ngat), .B(G2963_1741_ngat), .Y(G2965_1805_gat) );
OR2XL U_g1606 (.A(G1804_1513_ngat), .B(G1803_1152_ngat), .Y(G1805_1806_gat) );
OR2XL U_g1607 (.A(G1555_1514_ngat), .B(G1554_1153_ngat), .Y(G1556_1807_gat) );
OR2XL U_g1608 (.A(G2972_1515_ngat), .B(G2971_1744_ngat), .Y(G2973_1808_gat) );
OR2XL U_g1609 (.A(G7496_1516_ngat), .B(G7495_1523_ngat), .Y(G7598_1809_gat) );
OR2XL U_g1610 (.A(G1572_1517_ngat), .B(G1571_1156_ngat), .Y(G1573_1810_gat) );
OR2XL U_g1611 (.A(G1821_1518_ngat), .B(G1820_1157_ngat), .Y(G1822_1811_gat) );
OR2XL U_g1612 (.A(G1849_1521_ngat), .B(G1848_1160_ngat), .Y(G1850_1812_gat) );
OR2XL U_g1613 (.A(G1686_1522_ngat), .B(G1685_1163_ngat), .Y(G1687_1813_gat) );
OR2XL U_g1614 (.A(G3017_1524_ngat), .B(G3016_1745_ngat), .Y(G3018_1814_gat) );
OR2XL U_g1615 (.A(G4548_1525_ngat), .B(G4547_1532_ngat), .Y(G4549_1815_gat) );
OR2XL U_g1616 (.A(G2981_1526_ngat), .B(G2980_1748_ngat), .Y(G2982_1816_gat) );
OR2XL U_g1617 (.A(G1597_1527_ngat), .B(G1596_1168_ngat), .Y(G1598_1817_gat) );
OR2XL U_g1618 (.A(G1858_1528_ngat), .B(G1857_1169_ngat), .Y(G1859_1818_gat) );
OR2XL U_g1619 (.A(G1868_1529_ngat), .B(G1867_1170_ngat), .Y(G1869_1819_gat) );
OR2XL U_g1620 (.A(G1608_1530_ngat), .B(G1607_1171_ngat), .Y(G1609_1820_gat) );
OR2XL U_g1621 (.A(G2991_1531_ngat), .B(G2990_1579_ngat), .Y(G2992_1821_gat) );
OR2XL U_g1622 (.A(G4539_1533_ngat), .B(G4538_1540_ngat), .Y(G4540_1822_gat) );
OR2XL U_g1623 (.A(G3000_1534_ngat), .B(G2999_1578_ngat), .Y(G3001_1823_gat) );
OR2XL U_g1624 (.A(G1629_1535_ngat), .B(G1628_1176_ngat), .Y(G1630_1824_gat) );
OR2XL U_g1625 (.A(G1884_1536_ngat), .B(G1883_1177_ngat), .Y(G1885_1825_gat) );
OR2XL U_g1626 (.A(G1902_1537_ngat), .B(G1901_1178_ngat), .Y(G1903_1826_gat) );
OR2XL U_g1627 (.A(G1654_1538_ngat), .B(G1653_1179_ngat), .Y(G1655_1827_gat) );
OR2XL U_g1628 (.A(G3008_1539_ngat), .B(G3007_1575_ngat), .Y(G3009_1828_gat) );
OR2XL U_g1629 (.A(G1694_1542_ngat), .B(G1693_1184_ngat), .Y(G1695_1829_gat) );
OR2XL U_g1630 (.A(G4530_1185_ngat), .B(G4529_1545_ngat), .Y(G4531_1830_gat) );
OR2XL U_g1631 (.A(G3020_1543_ngat), .B(G3019_1581_ngat), .Y(G3021_1831_gat) );
OR2XL U_g1632 (.A(G1920_1544_ngat), .B(G1919_1188_ngat), .Y(G1921_1832_gat) );
INVXL U_g1633 (.A(G6832_1546_gat), .Y(G6836_1833_gat) );
INVXL U_g1634 (.A(G4932_1547_gat), .Y(G4936_1834_gat) );
INVXL U_g1635 (.A(G4973_1548_gat), .Y(G4977_1835_gat) );
OR2XL U_g1636 (.A(G906_1554_ngat), .B(G912_1550_ngat), .Y(G957_1836_gat) );
INVXL U_g1637 (.A(G4942_1551_gat), .Y(G4946_1837_gat) );
OR2XL U_g1638 (.A(G1112_1553_ngat), .B(G1121_1552_ngat), .Y(G1176_1838_gat) );
OR2XL U_g1639 (.A(G3521_1557_ngat), .B(G3520_1564_ngat), .Y(G3522_1839_gat) );
OR2XL U_g1640 (.A(G3175_1558_ngat), .B(G3174_1738_ngat), .Y(G3176_1840_gat) );
OR2XL U_g1641 (.A(G791_1559_ngat), .B(G790_1208_ngat), .Y(G792_1841_gat) );
OR2XL U_g1642 (.A(G1025_1560_ngat), .B(G1024_1209_ngat), .Y(G1026_1842_gat) );
OR2XL U_g1643 (.A(G1037_1561_ngat), .B(G1036_1210_ngat), .Y(G1038_1843_gat) );
OR2XL U_g1644 (.A(G804_1562_ngat), .B(G803_1211_ngat), .Y(G805_1844_gat) );
OR2XL U_g1645 (.A(G3185_1563_ngat), .B(G3184_1729_ngat), .Y(G3186_1845_gat) );
OR2XL U_g1646 (.A(G1073_1565_ngat), .B(G1072_1214_ngat), .Y(G1074_1846_gat) );
OR2XL U_g1647 (.A(G3202_1566_ngat), .B(G3201_1733_ngat), .Y(G3203_1847_gat) );
OR2XL U_g1648 (.A(G3512_1616_ngat), .B(G3511_1567_ngat), .Y(G3513_1848_gat) );
OR2XL U_g1649 (.A(G852_1568_ngat), .B(G851_1217_ngat), .Y(G853_1849_gat) );
OR2XL U_g1650 (.A(G894_1570_ngat), .B(G893_1220_ngat), .Y(G895_1850_gat) );
OR2XL U_g1651 (.A(G3503_1221_ngat), .B(G3502_1573_ngat), .Y(G3504_1851_gat) );
OR2XL U_g1652 (.A(G3214_1571_ngat), .B(G3213_1735_ngat), .Y(G3215_1852_gat) );
OR2XL U_g1653 (.A(G1092_1572_ngat), .B(G1091_1224_ngat), .Y(G1093_1853_gat) );
OR2XL U_g1654 (.A(G4225_1225_ngat), .B(G4224_1574_ngat), .Y(G4226_1854_gat) );
OR2XL U_g1655 (.A(G4234_1577_ngat), .B(G4233_1576_ngat), .Y(G4235_1855_gat) );
OR2XL U_g1656 (.A(G4243_1747_ngat), .B(G4242_1580_ngat), .Y(G4244_1856_gat) );
OR2XL U_g1657 (.A(G1262_1234_ngat), .B(G1261_1582_ngat), .Y(G1263_1857_gat) );
OR2XL U_g1658 (.A(G1271_1584_ngat), .B(G1270_1583_ngat), .Y(G1272_1858_gat) );
OR2XL U_g1659 (.A(G1280_1751_ngat), .B(G1279_1585_ngat), .Y(G1281_1859_gat) );
OR2XL U_g1660 (.A(G7279_1595_ngat), .B(G7276_1247_ngat), .Y(G7281_1860_gat) );
OR2XL U_g1661 (.A(G7423_1687_ngat), .B(G7420_1249_ngat), .Y(G4350_1861_gat) );
OR2XL U_g1662 (.A(G6795_1591_ngat), .B(G6792_1252_ngat), .Y(G6797_1862_gat) );
OR2XL U_g1663 (.A(G6796_1590_ngat), .B(G6789_1253_ngat), .Y(G6798_1863_gat) );
OR2XL U_g1664 (.A(G7383_1685_ngat), .B(G7380_1257_ngat), .Y(G4306_1864_gat) );
OR2XL U_g1665 (.A(G7280_1586_ngat), .B(G7273_1258_ngat), .Y(G7282_1865_gat) );
OR2XL U_g1666 (.A(G6805_1624_ngat), .B(G6802_1261_ngat), .Y(G6807_1866_gat) );
OR2XL U_g1667 (.A(G7375_1682_ngat), .B(G7372_1263_ngat), .Y(G4298_1867_gat) );
OR2XL U_g1668 (.A(G7289_1628_ngat), .B(G7286_1264_ngat), .Y(G7291_1868_gat) );
OR2XL U_g1669 (.A(G6743_1693_ngat), .B(G6740_1265_ngat), .Y(G3543_1869_gat) );
OR2XL U_g1670 (.A(G6477_1639_ngat), .B(G6474_1269_ngat), .Y(G3091_1870_gat) );
OR2XL U_g1671 (.A(G6509_1649_ngat), .B(G6506_1272_ngat), .Y(G3120_1871_gat) );
OR2XL U_g1672 (.A(G7211_1609_ngat), .B(G7208_978_ngat), .Y(G4178_1872_gat) );
OR2XL U_g1673 (.A(G6727_1611_ngat), .B(G6724_979_ngat), .Y(G3525_1873_gat) );
OR2XL U_g1674 (.A(G826_1614_ngat), .B(G825_1279_ngat), .Y(G827_1874_gat) );
OR2XL U_g1675 (.A(G1054_1615_ngat), .B(G1053_1280_ngat), .Y(G1055_1875_gat) );
OR2XL U_g1676 (.A(G3194_1617_ngat), .B(G3193_1731_ngat), .Y(G3195_1876_gat) );
OR2XL U_g1677 (.A(G7391_1662_ngat), .B(G7388_1283_ngat), .Y(G4315_1877_gat) );
OR2XL U_g1678 (.A(G6788_1719_ngat), .B(G6781_1286_ngat), .Y(G3567_1878_gat) );
OR2XL U_g1679 (.A(G6806_1598_ngat), .B(G6799_1289_ngat), .Y(G6808_1879_gat) );
OR2XL U_g1680 (.A(G7367_1681_ngat), .B(G7364_1292_ngat), .Y(G4289_1880_gat) );
OR2XL U_g1681 (.A(G7290_1600_ngat), .B(G7283_1294_ngat), .Y(G7292_1881_gat) );
OR2XL U_g1682 (.A(G6735_1634_ngat), .B(G6732_1295_ngat), .Y(G3534_1882_gat) );
OR2XL U_g1683 (.A(G6493_1647_ngat), .B(G6490_1299_ngat), .Y(G3108_1883_gat) );
OR2XL U_g1684 (.A(G7219_1638_ngat), .B(G7216_1300_ngat), .Y(G4187_1884_gat) );
OR2XL U_g1685 (.A(G6736_1629_ngat), .B(G6729_1301_ngat), .Y(G3535_1885_gat) );
OR2XL U_g1686 (.A(G6485_1678_ngat), .B(G6482_1304_ngat), .Y(G3100_1886_gat) );
OR2XL U_g1687 (.A(G7220_1633_ngat), .B(G7213_1306_ngat), .Y(G4188_1887_gat) );
OR2XL U_g1688 (.A(G6478_1604_ngat), .B(G6471_1307_ngat), .Y(G3092_1888_gat) );
OR2XL U_g1689 (.A(G7573_1643_ngat), .B(G7570_1308_ngat), .Y(G4593_1889_gat) );
OR2XL U_g1690 (.A(G7574_1640_ngat), .B(G7567_1310_ngat), .Y(G4594_1890_gat) );
OR2XL U_g1691 (.A(G7581_1677_ngat), .B(G7578_1312_ngat), .Y(G7583_1891_gat) );
OR2XL U_g1692 (.A(G6494_1632_ngat), .B(G6487_1313_ngat), .Y(G3109_1892_gat) );
OR2XL U_g1693 (.A(G7565_1679_ngat), .B(G7562_1314_ngat), .Y(G4584_1893_gat) );
OR2XL U_g1694 (.A(G6510_1607_ngat), .B(G6503_1315_ngat), .Y(G3121_1894_gat) );
OR2XL U_g1695 (.A(G7522_1660_ngat), .B(G7515_1317_ngat), .Y(G4562_1895_gat) );
OR2XL U_g1696 (.A(G7529_1661_ngat), .B(G7526_1320_ngat), .Y(G4570_1896_gat) );
OR2XL U_g1697 (.A(G7521_1652_ngat), .B(G7518_1322_ngat), .Y(G4561_1897_gat) );
OR2XL U_g1698 (.A(G7530_1657_ngat), .B(G7523_1323_ngat), .Y(G4571_1898_gat) );
OR2XL U_g1699 (.A(G7392_1618_ngat), .B(G7385_1324_ngat), .Y(G4316_1899_gat) );
OR2XL U_g1700 (.A(G4553_1663_ngat), .B(G4552_1664_ngat), .Y(G4554_1900_gat) );
OR2XL U_g1701 (.A(G6762_1689_ngat), .B(G6755_1328_ngat), .Y(G6764_1901_gat) );
OR2XL U_g1702 (.A(G7248_1668_ngat), .B(G7247_1691_ngat), .Y(G7337_1902_gat) );
OR2XL U_g1703 (.A(G6445_1670_ngat), .B(G6442_1006_ngat), .Y(G3050_1903_gat) );
OR2XL U_g1704 (.A(G7592_1674_ngat), .B(G7585_1334_ngat), .Y(G7594_1904_gat) );
OR2XL U_g1705 (.A(G7591_1671_ngat), .B(G7588_1336_ngat), .Y(G7593_1905_gat) );
OR2XL U_g1706 (.A(G7582_1646_ngat), .B(G7575_1338_ngat), .Y(G7584_1906_gat) );
OR2XL U_g1707 (.A(G6486_1637_ngat), .B(G6479_1339_ngat), .Y(G3101_1907_gat) );
OR2XL U_g1708 (.A(G7566_1648_ngat), .B(G7559_1340_ngat), .Y(G4585_1908_gat) );
OR2XL U_g1709 (.A(G7557_1651_ngat), .B(G7554_1011_ngat), .Y(G4575_1909_gat) );
OR2XL U_g1710 (.A(G7548_1683_ngat), .B(G7541_1342_ngat), .Y(G7550_1910_gat) );
OR2XL U_g1711 (.A(G7368_1627_ngat), .B(G7361_1343_ngat), .Y(G4290_1911_gat) );
OR2XL U_g1712 (.A(G7376_1599_ngat), .B(G7369_1344_ngat), .Y(G4299_1912_gat) );
OR2XL U_g1713 (.A(G7547_1680_ngat), .B(G7544_1345_ngat), .Y(G7549_1913_gat) );
OR2XL U_g1714 (.A(G7538_1686_ngat), .B(G7531_1346_ngat), .Y(G7540_1914_gat) );
OR2XL U_g1715 (.A(G7384_1594_ngat), .B(G7377_1347_ngat), .Y(G4307_1915_gat) );
OR2XL U_g1716 (.A(G7537_1684_ngat), .B(G7534_1348_ngat), .Y(G7539_1916_gat) );
OR2XL U_g1717 (.A(G7424_1587_ngat), .B(G7417_1349_ngat), .Y(G4351_1917_gat) );
OR2XL U_g1718 (.A(G6761_1666_ngat), .B(G6758_1351_ngat), .Y(G6763_1918_gat) );
OR2XL U_g1719 (.A(G6453_1673_ngat), .B(G6450_1017_ngat), .Y(G3060_1919_gat) );
OR2XL U_g1720 (.A(G6469_1642_ngat), .B(G6466_1019_ngat), .Y(G3080_1920_gat) );
OR2XL U_g1721 (.A(G7228_1606_ngat), .B(G7221_1020_ngat), .Y(G4197_1921_gat) );
OR2XL U_g1722 (.A(G6744_1601_ngat), .B(G6737_1360_ngat), .Y(G3544_1922_gat) );
OR2XL U_g1723 (.A(G4202_1362_ngat), .B(G4201_1695_ngat), .Y(G4203_1923_gat) );
OR2XL U_g1724 (.A(G6771_1697_ngat), .B(G6768_1023_ngat), .Y(G3548_1924_gat) );
INVXL U_g1725 (.A(G3223_1698_gat), .Y(G3227_1925_gat) );
OR2XL U_g1726 (.A(G4976_829_ngat), .B(G4973_1548_ngat), .Y(G4978_1926_gat) );
OR2XL U_g1727 (.A(G1157_1699_ngat), .B(G1156_1368_ngat), .Y(G1158_1927_gat) );
OR2XL U_g1728 (.A(G1153_1700_ngat), .B(G1152_1369_ngat), .Y(G1154_1928_gat) );
OR2XL U_g1729 (.A(G4935_722_ngat), .B(G4932_1547_ngat), .Y(G4937_1929_gat) );
OR2XL U_g1730 (.A(G6501_1645_ngat), .B(G6498_1032_ngat), .Y(G3117_1930_gat) );
OR2XL U_g1731 (.A(G7238_1708_ngat), .B(G7237_1701_ngat), .Y(G7340_1931_gat) );
OR2XL U_g1732 (.A(G6751_1705_ngat), .B(G6748_1373_ngat), .Y(G6753_1932_gat) );
OR2XL U_g1733 (.A(G6752_1702_ngat), .B(G6745_1376_ngat), .Y(G6754_1933_gat) );
OR2XL U_g1734 (.A(G6461_1676_ngat), .B(G6458_1036_ngat), .Y(G3069_1934_gat) );
OR2XL U_g1735 (.A(G6779_1713_ngat), .B(G6776_1384_ngat), .Y(G3557_1935_gat) );
OR2XL U_g1736 (.A(G7415_1659_ngat), .B(G7412_1039_ngat), .Y(G4342_1936_gat) );
OR2XL U_g1737 (.A(G4211_1716_ngat), .B(G4210_1712_ngat), .Y(G4212_1937_gat) );
OR2XL U_g1738 (.A(G6780_1711_ngat), .B(G6773_1388_ngat), .Y(G3558_1938_gat) );
OR2XL U_g1739 (.A(G7407_1654_ngat), .B(G7404_1042_ngat), .Y(G4334_1939_gat) );
OR2XL U_g1740 (.A(G6787_1621_ngat), .B(G6784_1396_ngat), .Y(G3566_1940_gat) );
OR2XL U_g1741 (.A(G7399_1656_ngat), .B(G7396_1045_ngat), .Y(G4325_1941_gat) );
OR2XL U_g1742 (.A(G7271_1620_ngat), .B(G7268_1046_ngat), .Y(G4219_1942_gat) );
OR2XL U_g1743 (.A(G7432_1724_ngat), .B(G7425_1047_ngat), .Y(G4354_1943_gat) );
BUFX20 U_g1744 (.A(G2724_1722_gat), .Y(G6261_1944_gat) );
OR2XL U_g1745 (.A(G5935_1402_ngat), .B(G5932_1726_ngat), .Y(G2470_1945_gat) );
INVXL U_g1746 (.A(G6173_1723_gat), .Y(G6179_1946_gat) );
OR2XL U_g1747 (.A(G6055_1403_ngat), .B(G6052_1725_ngat), .Y(G2740_1947_gat) );
INVXL U_g1748 (.A(G6052_1725_gat), .Y(G6056_1948_gat) );
INVXL U_g1749 (.A(G5932_1726_gat), .Y(G5936_1949_gat) );
OR2XL U_g1750 (.A(G1239_1734_ngat), .B(G1238_1727_ngat), .Y(G1240_1950_gat) );
OR2XL U_g1751 (.A(G1257_1737_ngat), .B(G1256_1728_ngat), .Y(G1258_1951_gat) );
OR2XL U_g1752 (.A(G1248_1730_ngat), .B(G1247_1732_ngat), .Y(G1249_1952_gat) );
INVXL U_g1753 (.A(G5380_1736_gat), .Y(G5384_1953_gat) );
OR2XL U_g1754 (.A(G7336_1739_ngat), .B(G7335_1742_ngat), .Y(G7353_1954_gat) );
OR2XL U_g1755 (.A(G7326_1743_ngat), .B(G7325_1746_ngat), .Y(G7356_1955_gat) );
OR2XL U_g1756 (.A(G5348_1749_ngat), .B(G5347_1750_ngat), .Y(G5362_1956_gat) );
OR2XL U_g1757 (.A(G5358_1752_ngat), .B(G5357_1753_ngat), .Y(G5359_1957_gat) );
OR2XL U_g1758 (.A(G1234_1760_ngat), .B(G1233_1754_ngat), .Y(G1235_1958_gat) );
OR2XL U_g1759 (.A(G1225_1755_ngat), .B(G1224_1756_ngat), .Y(G1226_1959_gat) );
OR2XL U_g1760 (.A(G1216_1757_ngat), .B(G1215_1758_ngat), .Y(G1217_1960_gat) );
INVXL U_g1761 (.A(G5372_1759_gat), .Y(G5376_1961_gat) );
OR2XL U_g1762 (.A(G3220_1761_ngat), .B(G3227_1925_ngat), .Y(G3244_1962_gat) );
OR2XL U_g1763 (.A(G3844_1762_ngat), .B(G3843_1463_ngat), .Y(G3845_1963_gat) );
OR2XL U_g1764 (.A(G3282_1763_ngat), .B(G3281_1464_ngat), .Y(G3283_1964_gat) );
OR2XL U_g1765 (.A(G3294_1764_ngat), .B(G3293_1465_ngat), .Y(G3295_1965_gat) );
OR2XL U_g1766 (.A(G3855_1765_ngat), .B(G3854_1466_ngat), .Y(G3856_1966_gat) );
OR2XL U_g1767 (.A(G3313_1766_ngat), .B(G3312_1467_ngat), .Y(G3314_1967_gat) );
OR2XL U_g1768 (.A(G3873_1767_ngat), .B(G3872_1468_ngat), .Y(G3874_1968_gat) );
OR2XL U_g1769 (.A(G3988_1770_ngat), .B(G3987_1472_ngat), .Y(G3989_1969_gat) );
OR2XL U_g1770 (.A(G3343_1771_ngat), .B(G3342_1473_ngat), .Y(G3344_1970_gat) );
OR2XL U_g1771 (.A(G3898_1772_ngat), .B(G3897_1475_ngat), .Y(G3899_1971_gat) );
OR2XL U_g1772 (.A(G3352_1773_ngat), .B(G3351_1476_ngat), .Y(G3353_1972_gat) );
OR2XL U_g1773 (.A(G3364_1774_ngat), .B(G3363_1477_ngat), .Y(G3365_1973_gat) );
OR2XL U_g1774 (.A(G3910_1775_ngat), .B(G3909_1478_ngat), .Y(G3911_1974_gat) );
OR2XL U_g1775 (.A(G3931_1776_ngat), .B(G3930_1479_ngat), .Y(G3932_1975_gat) );
OR2XL U_g1776 (.A(G3380_1777_ngat), .B(G3379_1480_ngat), .Y(G3381_1976_gat) );
OR2XL U_g1777 (.A(G3956_1778_ngat), .B(G3955_1481_ngat), .Y(G3957_1977_gat) );
OR2XL U_g1778 (.A(G3398_1779_ngat), .B(G3397_1482_ngat), .Y(G3399_1978_gat) );
OR2XL U_g1779 (.A(G3416_1781_ngat), .B(G3415_1484_ngat), .Y(G3417_1979_gat) );
OR2XL U_g1780 (.A(G3996_1782_ngat), .B(G3995_1486_ngat), .Y(G3997_1980_gat) );
OR2XL U_g1781 (.A(G2588_1783_ngat), .B(G2587_1487_ngat), .Y(G2589_1981_gat) );
OR2XL U_g1782 (.A(G2342_1784_ngat), .B(G2341_1488_ngat), .Y(G2343_1982_gat) );
OR2XL U_g1783 (.A(G2353_1785_ngat), .B(G2352_1489_ngat), .Y(G2354_1983_gat) );
OR2XL U_g1784 (.A(G2599_1786_ngat), .B(G2598_1490_ngat), .Y(G2600_1984_gat) );
OR2XL U_g1785 (.A(G2617_1787_ngat), .B(G2616_1491_ngat), .Y(G2618_1985_gat) );
OR2XL U_g1786 (.A(G2371_1788_ngat), .B(G2370_1492_ngat), .Y(G2372_1986_gat) );
OR2XL U_g1787 (.A(G2733_1791_ngat), .B(G2732_1496_ngat), .Y(G2734_1987_gat) );
OR2XL U_g1788 (.A(G2399_1792_ngat), .B(G2398_1497_ngat), .Y(G2400_1988_gat) );
OR2XL U_g1789 (.A(G2408_1793_ngat), .B(G2407_1499_ngat), .Y(G2409_1989_gat) );
OR2XL U_g1790 (.A(G2642_1794_ngat), .B(G2641_1500_ngat), .Y(G2643_1990_gat) );
OR2XL U_g1791 (.A(G2654_1795_ngat), .B(G2653_1501_ngat), .Y(G2655_1991_gat) );
OR2XL U_g1792 (.A(G2419_1796_ngat), .B(G2418_1502_ngat), .Y(G2420_1992_gat) );
OR2XL U_g1793 (.A(G2435_1797_ngat), .B(G2434_1503_ngat), .Y(G2436_1993_gat) );
OR2XL U_g1794 (.A(G2675_1798_ngat), .B(G2674_1504_ngat), .Y(G2676_1994_gat) );
OR2XL U_g1795 (.A(G2700_1799_ngat), .B(G2699_1505_ngat), .Y(G2701_1995_gat) );
OR2XL U_g1796 (.A(G2453_1800_ngat), .B(G2452_1506_ngat), .Y(G2454_1996_gat) );
INVXL U_g1797 (.A(G7595_1801_gat), .Y(G7601_1997_gat) );
AND4XL U_g1798 (.A(G2956_1802_gat), .B(G2965_1805_gat), .C(G2973_1808_gat), .D(G3018_1814_gat), .Y(G3022_1998_gat) );
AND4XL U_g1799 (.A(G1546_1803_gat), .B(G1556_1807_gat), .C(G1573_1810_gat), .D(G1687_1813_gat), .Y(G1702_1999_gat) );
BUFX20 U_g1800 (.A(G1546_1803_gat), .Y(G5566_2000_gat) );
BUFX20 U_g1801 (.A(G1546_1803_gat), .Y(G5508_2001_gat) );
BUFX20 U_g1802 (.A(G1795_1804_gat), .Y(G5820_2002_gat) );
BUFX20 U_g1803 (.A(G1795_1804_gat), .Y(G5828_2003_gat) );
AND4XL U_g1804 (.A(G1795_1804_gat), .B(G1822_1811_gat), .C(G1850_1812_gat), .D(G1805_1806_gat), .Y(G1935_2004_gat) );
AND2XL U_g1805 (.A(G2970_872_gat), .B(G2956_1802_gat), .Y(G3025_2005_gat) );
AND2XL U_g1806 (.A(G1816_875_gat), .B(G1795_1804_gat), .Y(G1938_2006_gat) );
BUFX20 U_g1807 (.A(G1805_1806_gat), .Y(G5844_2007_gat) );
BUFX20 U_g1808 (.A(G1805_1806_gat), .Y(G5836_2008_gat) );
AND3XL U_g1809 (.A(G1805_1806_gat), .B(G1822_1811_gat), .C(G1850_1812_gat), .Y(G1944_2009_gat) );
AND2XL U_g1810 (.A(G1567_876_gat), .B(G1546_1803_gat), .Y(G1705_2010_gat) );
BUFX20 U_g1811 (.A(G1556_1807_gat), .Y(G5518_2011_gat) );
AND3XL U_g1812 (.A(G1556_1807_gat), .B(G1573_1810_gat), .C(G1687_1813_gat), .Y(G1711_2012_gat) );
BUFX20 U_g1813 (.A(G1556_1807_gat), .Y(G5576_2013_gat) );
AND2XL U_g1814 (.A(G1584_877_gat), .B(G1556_1807_gat), .Y(G1712_2014_gat) );
AND3XL U_g1815 (.A(G1584_877_gat), .B(G1546_1803_gat), .C(G1556_1807_gat), .Y(G1706_2015_gat) );
AND2XL U_g1816 (.A(G1584_877_gat), .B(G1556_1807_gat), .Y(G1709_2016_gat) );
AND3XL U_g1817 (.A(G1834_878_gat), .B(G1795_1804_gat), .C(G1805_1806_gat), .Y(G1939_2017_gat) );
AND2XL U_g1818 (.A(G1834_878_gat), .B(G1805_1806_gat), .Y(G1942_2018_gat) );
AND2XL U_g1819 (.A(G1834_878_gat), .B(G1805_1806_gat), .Y(G1945_2019_gat) );
AND3XL U_g1820 (.A(G2977_879_gat), .B(G2956_1802_gat), .C(G2965_1805_gat), .Y(G3026_2020_gat) );
INVXL U_g1821 (.A(G7598_1809_gat), .Y(G7602_2021_gat) );
AND2XL U_g1822 (.A(G1573_1810_gat), .B(G1687_1813_gat), .Y(G1749_2022_gat) );
BUFX20 U_g1823 (.A(G1573_1810_gat), .Y(G5498_2023_gat) );
BUFX20 U_g1824 (.A(G1573_1810_gat), .Y(G5556_2024_gat) );
BUFX20 U_g1825 (.A(G1822_1811_gat), .Y(G5860_2025_gat) );
BUFX20 U_g1826 (.A(G1822_1811_gat), .Y(G5852_2026_gat) );
AND2XL U_g1827 (.A(G1822_1811_gat), .B(G1850_1812_gat), .Y(G1948_2027_gat) );
AND3XL U_g1828 (.A(G1556_1807_gat), .B(G1590_882_gat), .C(G1573_1810_gat), .Y(G1710_2028_gat) );
AND4XL U_g1829 (.A(G1556_1807_gat), .B(G1590_882_gat), .C(G1546_1803_gat), .D(G1573_1810_gat), .Y(G1707_2029_gat) );
AND3XL U_g1830 (.A(G1556_1807_gat), .B(G1590_882_gat), .C(G1573_1810_gat), .Y(G1713_2030_gat) );
AND2XL U_g1831 (.A(G1590_882_gat), .B(G1573_1810_gat), .Y(G1714_2031_gat) );
AND4XL U_g1832 (.A(G1805_1806_gat), .B(G1841_883_gat), .C(G1795_1804_gat), .D(G1822_1811_gat), .Y(G1940_2032_gat) );
AND3XL U_g1833 (.A(G1805_1806_gat), .B(G1822_1811_gat), .C(G1841_883_gat), .Y(G1946_2033_gat) );
AND3XL U_g1834 (.A(G1805_1806_gat), .B(G1841_883_gat), .C(G1822_1811_gat), .Y(G1943_2034_gat) );
AND2XL U_g1835 (.A(G1841_883_gat), .B(G1822_1811_gat), .Y(G1947_2035_gat) );
AND2XL U_g1836 (.A(G1841_883_gat), .B(G1822_1811_gat), .Y(G1949_2036_gat) );
INVXL U_g1837 (.A(G1850_1812_gat), .Y(G1856_2037_gat) );
BUFX20 U_g1838 (.A(G1687_1813_gat), .Y(G5546_2038_gat) );
BUFX20 U_g1839 (.A(G1687_1813_gat), .Y(G5488_2039_gat) );
AND4XL U_g1840 (.A(G2965_1805_gat), .B(G2979_886_gat), .C(G2956_1802_gat), .D(G2973_1808_gat), .Y(G3027_2040_gat) );
BUFX20 U_g1841 (.A(G4549_1815_gat), .Y(G4602_2041_gat) );
BUFX20 U_g1842 (.A(G4549_1815_gat), .Y(G4598_2042_gat) );
AND5XL U_g1843 (.A(G2982_1816_gat), .B(G2992_1821_gat), .C(G3001_1823_gat), .D(G3009_1828_gat), .E(G3021_1831_gat), .Y(G3029_2043_gat) );
BUFX20 U_g1844 (.A(G1598_1817_gat), .Y(G5722_2044_gat) );
BUFX20 U_g1845 (.A(G1598_1817_gat), .Y(G5634_2045_gat) );
AND5XL U_g1846 (.A(G1598_1817_gat), .B(G1609_1820_gat), .C(G1630_1824_gat), .D(G1655_1827_gat), .E(G1695_1829_gat), .Y(G1718_2046_gat) );
AND5XL U_g1847 (.A(G1903_1826_gat), .B(G1859_1818_gat), .C(G1885_1825_gat), .D(G1921_1832_gat), .E(G1869_1819_gat), .Y(G1950_2047_gat) );
BUFX20 U_g1848 (.A(G1859_1818_gat), .Y(G4724_2048_gat) );
AND2XL U_g1849 (.A(G1624_894_gat), .B(G1598_1817_gat), .Y(G1722_2049_gat) );
AND2XL U_g1850 (.A(G1880_895_gat), .B(G1859_1818_gat), .Y(G1953_2050_gat) );
BUFX20 U_g1851 (.A(G1869_1819_gat), .Y(G4732_2051_gat) );
BUFX20 U_g1852 (.A(G1609_1820_gat), .Y(G5664_2052_gat) );
AND4XL U_g1853 (.A(G1655_1827_gat), .B(G1609_1820_gat), .C(G1630_1824_gat), .D(G1695_1829_gat), .Y(G1736_2053_gat) );
BUFX20 U_g1854 (.A(G1609_1820_gat), .Y(G5654_2054_gat) );
AND2XL U_g1855 (.A(G2998_896_gat), .B(G2982_1816_gat), .Y(G3030_2055_gat) );
AND2XL U_g1856 (.A(G1647_899_gat), .B(G1609_1820_gat), .Y(G1737_2056_gat) );
AND2XL U_g1857 (.A(G1647_899_gat), .B(G1609_1820_gat), .Y(G1733_2057_gat) );
AND3XL U_g1858 (.A(G1647_899_gat), .B(G1598_1817_gat), .C(G1609_1820_gat), .Y(G1723_2058_gat) );
AND2XL U_g1859 (.A(G1897_900_gat), .B(G1869_1819_gat), .Y(G1960_2059_gat) );
AND3XL U_g1860 (.A(G1897_900_gat), .B(G1859_1818_gat), .C(G1869_1819_gat), .Y(G1954_2060_gat) );
AND3XL U_g1861 (.A(G3006_901_gat), .B(G2982_1816_gat), .C(G2992_1821_gat), .Y(G3031_2061_gat) );
INVXL U_g1862 (.A(G4540_1822_gat), .Y(G4544_2062_gat) );
BUFX20 U_g1863 (.A(G1630_1824_gat), .Y(G5732_2063_gat) );
BUFX20 U_g1864 (.A(G1630_1824_gat), .Y(G5644_2064_gat) );
AND3XL U_g1865 (.A(G1655_1827_gat), .B(G1630_1824_gat), .C(G1695_1829_gat), .Y(G1742_2065_gat) );
BUFX20 U_g1866 (.A(G1885_1825_gat), .Y(G4740_2066_gat) );
AND3XL U_g1867 (.A(G1609_1820_gat), .B(G1669_904_gat), .C(G1630_1824_gat), .Y(G1738_2067_gat) );
AND3XL U_g1868 (.A(G1609_1820_gat), .B(G1669_904_gat), .C(G1630_1824_gat), .Y(G1734_2068_gat) );
AND4XL U_g1869 (.A(G1609_1820_gat), .B(G1669_904_gat), .C(G1598_1817_gat), .D(G1630_1824_gat), .Y(G1724_2069_gat) );
AND2XL U_g1870 (.A(G1669_904_gat), .B(G1630_1824_gat), .Y(G1743_2070_gat) );
AND2XL U_g1871 (.A(G1669_904_gat), .B(G1630_1824_gat), .Y(G1740_2071_gat) );
AND3XL U_g1872 (.A(G1869_1819_gat), .B(G1914_905_gat), .C(G1885_1825_gat), .Y(G1961_2072_gat) );
AND4XL U_g1873 (.A(G1869_1819_gat), .B(G1914_905_gat), .C(G1859_1818_gat), .D(G1885_1825_gat), .Y(G1955_2073_gat) );
AND2XL U_g1874 (.A(G1885_1825_gat), .B(G1914_905_gat), .Y(G1965_2074_gat) );
BUFX20 U_g1875 (.A(G1903_1826_gat), .Y(G4748_2075_gat) );
BUFX20 U_g1876 (.A(G1655_1827_gat), .Y(G5624_2076_gat) );
BUFX20 U_g1877 (.A(G1655_1827_gat), .Y(G5712_2077_gat) );
AND2XL U_g1878 (.A(G1655_1827_gat), .B(G1695_1829_gat), .Y(G1750_2078_gat) );
AND4XL U_g1879 (.A(G2992_1821_gat), .B(G3013_906_gat), .C(G2982_1816_gat), .D(G3001_1823_gat), .Y(G3032_2079_gat) );
AND4XL U_g1880 (.A(G1609_1820_gat), .B(G1677_909_gat), .C(G1630_1824_gat), .D(G1655_1827_gat), .Y(G1735_2080_gat) );
AND5XL U_g1881 (.A(G1609_1820_gat), .B(G1677_909_gat), .C(G1598_1817_gat), .D(G1630_1824_gat), .E(G1655_1827_gat), .Y(G1725_2081_gat) );
AND4XL U_g1882 (.A(G1609_1820_gat), .B(G1677_909_gat), .C(G1630_1824_gat), .D(G1655_1827_gat), .Y(G1739_2082_gat) );
AND3XL U_g1883 (.A(G1677_909_gat), .B(G1630_1824_gat), .C(G1655_1827_gat), .Y(G1741_2083_gat) );
AND2XL U_g1884 (.A(G1677_909_gat), .B(G1655_1827_gat), .Y(G1745_2084_gat) );
AND3XL U_g1885 (.A(G1677_909_gat), .B(G1630_1824_gat), .C(G1655_1827_gat), .Y(G1744_2085_gat) );
AND4XL U_g1886 (.A(G1869_1819_gat), .B(G1929_910_gat), .C(G1885_1825_gat), .D(G1903_1826_gat), .Y(G1962_2086_gat) );
AND5XL U_g1887 (.A(G1869_1819_gat), .B(G1929_910_gat), .C(G1859_1818_gat), .D(G1885_1825_gat), .E(G1903_1826_gat), .Y(G1956_2087_gat) );
AND2XL U_g1888 (.A(G1929_910_gat), .B(G1903_1826_gat), .Y(G1969_2088_gat) );
AND3XL U_g1889 (.A(G1929_910_gat), .B(G1885_1825_gat), .C(G1903_1826_gat), .Y(G1966_2089_gat) );
BUFX20 U_g1890 (.A(G1695_1829_gat), .Y(G5702_2090_gat) );
BUFX20 U_g1891 (.A(G1695_1829_gat), .Y(G5614_2091_gat) );
AND5XL U_g1892 (.A(G2992_1821_gat), .B(G3015_912_gat), .C(G2982_1816_gat), .D(G3001_1823_gat), .E(G3009_1828_gat), .Y(G3033_2092_gat) );
INVXL U_g1893 (.A(G4531_1830_gat), .Y(G4535_2093_gat) );
BUFX20 U_g1894 (.A(G1921_1832_gat), .Y(G4716_2094_gat) );
BUFX20 U_g1895 (.A(G3522_1839_gat), .Y(G3575_2095_gat) );
BUFX20 U_g1896 (.A(G3522_1839_gat), .Y(G3571_2096_gat) );
AND5XL U_g1897 (.A(G3176_1840_gat), .B(G3186_1845_gat), .C(G3195_1876_gat), .D(G3203_1847_gat), .E(G3215_1852_gat), .Y(G3228_2097_gat) );
BUFX20 U_g1898 (.A(G792_1841_gat), .Y(G5152_2098_gat) );
BUFX20 U_g1899 (.A(G792_1841_gat), .Y(G5064_2099_gat) );
AND5XL U_g1900 (.A(G792_1841_gat), .B(G805_1844_gat), .C(G827_1874_gat), .D(G853_1849_gat), .E(G895_1850_gat), .Y(G920_2100_gat) );
AND5XL U_g1901 (.A(G1074_1846_gat), .B(G1026_1842_gat), .C(G1055_1875_gat), .D(G1093_1853_gat), .E(G1038_1843_gat), .Y(G1122_2101_gat) );
BUFX20 U_g1902 (.A(G1026_1842_gat), .Y(G4764_2102_gat) );
AND2XL U_g1903 (.A(G821_929_gat), .B(G792_1841_gat), .Y(G925_2103_gat) );
AND2XL U_g1904 (.A(G1050_930_gat), .B(G1026_1842_gat), .Y(G1125_2104_gat) );
BUFX20 U_g1905 (.A(G1038_1843_gat), .Y(G4772_2105_gat) );
BUFX20 U_g1906 (.A(G805_1844_gat), .Y(G5094_2106_gat) );
AND4XL U_g1907 (.A(G853_1849_gat), .B(G805_1844_gat), .C(G827_1874_gat), .D(G895_1850_gat), .Y(G940_2107_gat) );
BUFX20 U_g1908 (.A(G805_1844_gat), .Y(G5084_2108_gat) );
AND2XL U_g1909 (.A(G3192_931_gat), .B(G3176_1840_gat), .Y(G3231_2109_gat) );
AND3XL U_g1910 (.A(G805_1844_gat), .B(G868_934_gat), .C(G827_1874_gat), .Y(G942_2110_gat) );
AND3XL U_g1911 (.A(G805_1844_gat), .B(G868_934_gat), .C(G827_1874_gat), .Y(G938_2111_gat) );
AND4XL U_g1912 (.A(G805_1844_gat), .B(G868_934_gat), .C(G792_1841_gat), .D(G827_1874_gat), .Y(G927_2112_gat) );
AND2XL U_g1913 (.A(G868_934_gat), .B(G827_1874_gat), .Y(G947_2113_gat) );
AND2XL U_g1914 (.A(G868_934_gat), .B(G827_1874_gat), .Y(G944_2114_gat) );
AND3XL U_g1915 (.A(G1038_1843_gat), .B(G1086_935_gat), .C(G1055_1875_gat), .Y(G1133_2115_gat) );
AND4XL U_g1916 (.A(G1038_1843_gat), .B(G1086_935_gat), .C(G1026_1842_gat), .D(G1055_1875_gat), .Y(G1127_2116_gat) );
AND2XL U_g1917 (.A(G1055_1875_gat), .B(G1086_935_gat), .Y(G1137_2117_gat) );
BUFX20 U_g1918 (.A(G1074_1846_gat), .Y(G4788_2118_gat) );
AND4XL U_g1919 (.A(G3186_1845_gat), .B(G3207_936_gat), .C(G3176_1840_gat), .D(G3195_1876_gat), .Y(G3233_2119_gat) );
INVXL U_g1920 (.A(G3513_1848_gat), .Y(G3517_2120_gat) );
BUFX20 U_g1921 (.A(G853_1849_gat), .Y(G5054_2121_gat) );
AND3XL U_g1922 (.A(G853_1849_gat), .B(G827_1874_gat), .C(G895_1850_gat), .Y(G946_2122_gat) );
BUFX20 U_g1923 (.A(G853_1849_gat), .Y(G5142_2123_gat) );
AND2XL U_g1924 (.A(G853_1849_gat), .B(G895_1850_gat), .Y(G956_2124_gat) );
AND4XL U_g1925 (.A(G805_1844_gat), .B(G877_939_gat), .C(G827_1874_gat), .D(G853_1849_gat), .Y(G939_2125_gat) );
AND5XL U_g1926 (.A(G805_1844_gat), .B(G877_939_gat), .C(G792_1841_gat), .D(G827_1874_gat), .E(G853_1849_gat), .Y(G928_2126_gat) );
AND4XL U_g1927 (.A(G805_1844_gat), .B(G877_939_gat), .C(G827_1874_gat), .D(G853_1849_gat), .Y(G943_2127_gat) );
AND3XL U_g1928 (.A(G877_939_gat), .B(G827_1874_gat), .C(G853_1849_gat), .Y(G945_2128_gat) );
AND2XL U_g1929 (.A(G877_939_gat), .B(G853_1849_gat), .Y(G949_2129_gat) );
AND3XL U_g1930 (.A(G877_939_gat), .B(G827_1874_gat), .C(G853_1849_gat), .Y(G948_2130_gat) );
AND4XL U_g1931 (.A(G1038_1843_gat), .B(G1102_940_gat), .C(G1055_1875_gat), .D(G1074_1846_gat), .Y(G1134_2131_gat) );
AND5XL U_g1932 (.A(G1038_1843_gat), .B(G1102_940_gat), .C(G1026_1842_gat), .D(G1055_1875_gat), .E(G1074_1846_gat), .Y(G1128_2132_gat) );
AND2XL U_g1933 (.A(G1102_940_gat), .B(G1074_1846_gat), .Y(G1141_2133_gat) );
AND3XL U_g1934 (.A(G1102_940_gat), .B(G1055_1875_gat), .C(G1074_1846_gat), .Y(G1138_2134_gat) );
BUFX20 U_g1935 (.A(G895_1850_gat), .Y(G5132_2135_gat) );
BUFX20 U_g1936 (.A(G895_1850_gat), .Y(G5044_2136_gat) );
AND5XL U_g1937 (.A(G3186_1845_gat), .B(G3209_942_gat), .C(G3176_1840_gat), .D(G3195_1876_gat), .E(G3203_1847_gat), .Y(G3234_2137_gat) );
INVXL U_g1938 (.A(G3504_1851_gat), .Y(G3508_2138_gat) );
BUFX20 U_g1939 (.A(G1093_1853_gat), .Y(G4756_2139_gat) );
INVXL U_g1940 (.A(G4226_1854_gat), .Y(G4230_2140_gat) );
INVXL U_g1941 (.A(G4235_1855_gat), .Y(G4239_2141_gat) );
BUFX20 U_g1942 (.A(G4244_1856_gat), .Y(G4263_2142_gat) );
BUFX20 U_g1943 (.A(G4244_1856_gat), .Y(G4267_2143_gat) );
INVXL U_g1944 (.A(G1263_1857_gat), .Y(G1267_2144_gat) );
INVXL U_g1945 (.A(G1272_1858_gat), .Y(G1276_2145_gat) );
BUFX20 U_g1946 (.A(G1281_1859_gat), .Y(G1300_2146_gat) );
BUFX20 U_g1947 (.A(G1281_1859_gat), .Y(G1304_2147_gat) );
OR2XL U_g1948 (.A(G7282_1865_ngat), .B(G7281_1860_ngat), .Y(G7348_2148_gat) );
OR2XL U_g1949 (.A(G4351_1917_ngat), .B(G4350_1861_ngat), .Y(G4352_2149_gat) );
OR2XL U_g1950 (.A(G6798_1863_ngat), .B(G6797_1862_ngat), .Y(G6822_2150_gat) );
OR2XL U_g1951 (.A(G4307_1915_ngat), .B(G4306_1864_ngat), .Y(G4308_2151_gat) );
OR2XL U_g1952 (.A(G6808_1879_ngat), .B(G6807_1866_ngat), .Y(G6819_2152_gat) );
OR2XL U_g1953 (.A(G4299_1912_ngat), .B(G4298_1867_ngat), .Y(G4300_2153_gat) );
OR2XL U_g1954 (.A(G7292_1881_ngat), .B(G7291_1868_ngat), .Y(G7345_2154_gat) );
OR2XL U_g1955 (.A(G3544_1922_ngat), .B(G3543_1869_ngat), .Y(G3545_2155_gat) );
OR2XL U_g1956 (.A(G3092_1888_ngat), .B(G3091_1870_ngat), .Y(G3093_2156_gat) );
OR2XL U_g1957 (.A(G4197_1921_ngat), .B(G4196_1605_ngat), .Y(G4198_2157_gat) );
OR2XL U_g1958 (.A(G3121_1894_ngat), .B(G3120_1871_ngat), .Y(G3122_2158_gat) );
OR2XL U_g1959 (.A(G4179_1608_ngat), .B(G4178_1872_ngat), .Y(G4180_2159_gat) );
OR2XL U_g1960 (.A(G3526_1610_ngat), .B(G3525_1873_ngat), .Y(G3527_2160_gat) );
AND2XL U_g1961 (.A(G845_980_gat), .B(G805_1844_gat), .Y(G941_2161_gat) );
AND2XL U_g1962 (.A(G845_980_gat), .B(G805_1844_gat), .Y(G937_2162_gat) );
AND3XL U_g1963 (.A(G845_980_gat), .B(G792_1841_gat), .C(G805_1844_gat), .Y(G926_2163_gat) );
AND2XL U_g1964 (.A(G1068_981_gat), .B(G1038_1843_gat), .Y(G1132_2164_gat) );
AND3XL U_g1965 (.A(G1068_981_gat), .B(G1026_1842_gat), .C(G1038_1843_gat), .Y(G1126_2165_gat) );
BUFX20 U_g1966 (.A(G827_1874_gat), .Y(G5162_2166_gat) );
BUFX20 U_g1967 (.A(G827_1874_gat), .Y(G5074_2167_gat) );
BUFX20 U_g1968 (.A(G1055_1875_gat), .Y(G4780_2168_gat) );
AND3XL U_g1969 (.A(G3200_982_gat), .B(G3176_1840_gat), .C(G3186_1845_gat), .Y(G3232_2169_gat) );
OR2XL U_g1970 (.A(G4316_1899_ngat), .B(G4315_1877_ngat), .Y(G4317_2170_gat) );
OR2XL U_g1971 (.A(G4220_1619_ngat), .B(G4219_1942_ngat), .Y(G4221_2171_gat) );
OR2XL U_g1972 (.A(G3567_1878_ngat), .B(G3566_1940_ngat), .Y(G3568_2172_gat) );
OR2XL U_g1973 (.A(G4290_1911_ngat), .B(G4289_1880_ngat), .Y(G4291_2173_gat) );
OR2XL U_g1974 (.A(G3535_1885_ngat), .B(G3534_1882_ngat), .Y(G3536_2174_gat) );
OR2XL U_g1975 (.A(G3109_1892_ngat), .B(G3108_1883_ngat), .Y(G3110_2175_gat) );
OR2XL U_g1976 (.A(G4188_1887_ngat), .B(G4187_1884_ngat), .Y(G4189_2176_gat) );
OR2XL U_g1977 (.A(G3101_1907_ngat), .B(G3100_1886_ngat), .Y(G3102_2177_gat) );
OR2XL U_g1978 (.A(G4594_1890_ngat), .B(G4593_1889_ngat), .Y(G4595_2178_gat) );
OR2XL U_g1979 (.A(G3081_1641_ngat), .B(G3080_1920_ngat), .Y(G3082_2179_gat) );
OR2XL U_g1980 (.A(G3118_1644_ngat), .B(G3117_1930_ngat), .Y(G3119_2180_gat) );
OR2XL U_g1981 (.A(G7584_1906_ngat), .B(G7583_1891_ngat), .Y(G7614_2181_gat) );
OR2XL U_g1982 (.A(G4585_1908_ngat), .B(G4584_1893_ngat), .Y(G4586_2182_gat) );
OR2XL U_g1983 (.A(G4576_1650_ngat), .B(G4575_1909_ngat), .Y(G4577_2183_gat) );
OR2XL U_g1984 (.A(G4562_1895_ngat), .B(G4561_1897_ngat), .Y(G4563_2184_gat) );
OR2XL U_g1985 (.A(G4335_1653_ngat), .B(G4334_1939_ngat), .Y(G4336_2185_gat) );
OR2XL U_g1986 (.A(G4326_1655_ngat), .B(G4325_1941_ngat), .Y(G4327_2186_gat) );
OR2XL U_g1987 (.A(G4571_1898_ngat), .B(G4570_1896_ngat), .Y(G4572_2187_gat) );
OR2XL U_g1988 (.A(G4343_1658_ngat), .B(G4342_1936_ngat), .Y(G4344_2188_gat) );
INVXL U_g1989 (.A(G4554_1900_gat), .Y(G4558_2189_gat) );
OR2XL U_g1990 (.A(G6764_1901_ngat), .B(G6763_1918_ngat), .Y(G6809_2190_gat) );
INVXL U_g1991 (.A(G7337_1902_gat), .Y(G7343_2191_gat) );
OR2XL U_g1992 (.A(G3051_1669_ngat), .B(G3050_1903_ngat), .Y(G3052_2192_gat) );
OR2XL U_g1993 (.A(G7594_1904_ngat), .B(G7593_1905_ngat), .Y(G7611_2193_gat) );
OR2XL U_g1994 (.A(G3061_1672_ngat), .B(G3060_1919_ngat), .Y(G3062_2194_gat) );
OR2XL U_g1995 (.A(G3070_1675_ngat), .B(G3069_1934_ngat), .Y(G3071_2195_gat) );
OR2XL U_g1996 (.A(G7550_1910_ngat), .B(G7549_1913_ngat), .Y(G7603_2196_gat) );
OR2XL U_g1997 (.A(G7540_1914_ngat), .B(G7539_1916_ngat), .Y(G7606_2197_gat) );
INVXL U_g1998 (.A(G4203_1923_gat), .Y(G4207_2198_gat) );
OR2XL U_g1999 (.A(G3549_1696_ngat), .B(G3548_1924_ngat), .Y(G3550_2199_gat) );
OR2XL U_g2000 (.A(G4977_1835_ngat), .B(G4970_718_ngat), .Y(G4979_2200_gat) );
INVXL U_g2001 (.A(G1154_1928_gat), .Y(G1155_2201_gat) );
OR2XL U_g2002 (.A(G4936_1834_ngat), .B(G4929_564_ngat), .Y(G4938_2202_gat) );
INVXL U_g2003 (.A(G7340_1931_gat), .Y(G7344_2203_gat) );
OR2XL U_g2004 (.A(G6754_1933_ngat), .B(G6753_1932_ngat), .Y(G6812_2204_gat) );
OR2XL U_g2005 (.A(G3558_1938_ngat), .B(G3557_1935_ngat), .Y(G3559_2205_gat) );
INVXL U_g2006 (.A(G4212_1937_gat), .Y(G4216_2206_gat) );
OR2XL U_g2007 (.A(G4354_1943_ngat), .B(G4353_1720_ngat), .Y(G4355_2207_gat) );
INVXL U_g2008 (.A(G6261_1944_gat), .Y(G6267_2208_gat) );
OR2XL U_g2009 (.A(G5936_1949_ngat), .B(G5929_1048_ngat), .Y(G2471_2209_gat) );
OR2XL U_g2010 (.A(G6056_1948_ngat), .B(G6049_1049_ngat), .Y(G2741_2210_gat) );
INVXL U_g2011 (.A(G1240_1950_gat), .Y(G1244_2211_gat) );
BUFX20 U_g2012 (.A(G1258_1951_gat), .Y(G1296_2212_gat) );
BUFX20 U_g2013 (.A(G1258_1951_gat), .Y(G1292_2213_gat) );
INVXL U_g2014 (.A(G1249_1952_gat), .Y(G1253_2214_gat) );
INVXL U_g2015 (.A(G7353_1954_gat), .Y(G7359_2215_gat) );
INVXL U_g2016 (.A(G7356_1955_gat), .Y(G7360_2216_gat) );
INVXL U_g2017 (.A(G5362_1956_gat), .Y(G5366_2217_gat) );
INVXL U_g2018 (.A(G5359_1957_gat), .Y(G5365_2218_gat) );
BUFX20 U_g2019 (.A(G1235_1958_gat), .Y(G1288_2219_gat) );
BUFX20 U_g2020 (.A(G1235_1958_gat), .Y(G1284_2220_gat) );
INVXL U_g2021 (.A(G1226_1959_gat), .Y(G1230_2221_gat) );
INVXL U_g2022 (.A(G1217_1960_gat), .Y(G1221_2222_gat) );
AND2XL U_g2023 (.A(G3228_2097_gat), .B(G3216_1462_gat), .Y(G3249_2223_gat) );
AND4XL U_g2024 (.A(G3845_1963_gat), .B(G3856_1966_gat), .C(G3874_1968_gat), .D(G3989_1969_gat), .Y(G4004_2224_gat) );
BUFX20 U_g2025 (.A(G3845_1963_gat), .Y(G7026_2225_gat) );
BUFX20 U_g2026 (.A(G3845_1963_gat), .Y(G6968_2226_gat) );
BUFX20 U_g2027 (.A(G3283_1964_gat), .Y(G6642_2227_gat) );
BUFX20 U_g2028 (.A(G3283_1964_gat), .Y(G6650_2228_gat) );
AND4XL U_g2029 (.A(G3283_1964_gat), .B(G3314_1967_gat), .C(G3344_1970_gat), .D(G3295_1965_gat), .Y(G3431_2229_gat) );
AND2XL U_g2030 (.A(G3308_1109_gat), .B(G3283_1964_gat), .Y(G3434_2230_gat) );
AND2XL U_g2031 (.A(G3868_1110_gat), .B(G3845_1963_gat), .Y(G4007_2231_gat) );
BUFX20 U_g2032 (.A(G3295_1965_gat), .Y(G6666_2232_gat) );
BUFX20 U_g2033 (.A(G3295_1965_gat), .Y(G6658_2233_gat) );
AND3XL U_g2034 (.A(G3295_1965_gat), .B(G3314_1967_gat), .C(G3344_1970_gat), .Y(G3440_2234_gat) );
BUFX20 U_g2035 (.A(G3856_1966_gat), .Y(G6978_2235_gat) );
AND3XL U_g2036 (.A(G3856_1966_gat), .B(G3874_1968_gat), .C(G3989_1969_gat), .Y(G4013_2236_gat) );
BUFX20 U_g2037 (.A(G3856_1966_gat), .Y(G7036_2237_gat) );
AND3XL U_g2038 (.A(G3327_1111_gat), .B(G3283_1964_gat), .C(G3295_1965_gat), .Y(G3435_2238_gat) );
AND2XL U_g2039 (.A(G3327_1111_gat), .B(G3295_1965_gat), .Y(G3438_2239_gat) );
AND2XL U_g2040 (.A(G3327_1111_gat), .B(G3295_1965_gat), .Y(G3441_2240_gat) );
AND2XL U_g2041 (.A(G3885_1112_gat), .B(G3856_1966_gat), .Y(G4014_2241_gat) );
AND3XL U_g2042 (.A(G3885_1112_gat), .B(G3845_1963_gat), .C(G3856_1966_gat), .Y(G4008_2242_gat) );
AND2XL U_g2043 (.A(G3885_1112_gat), .B(G3856_1966_gat), .Y(G4011_2243_gat) );
BUFX20 U_g2044 (.A(G3314_1967_gat), .Y(G6682_2244_gat) );
BUFX20 U_g2045 (.A(G3314_1967_gat), .Y(G6674_2245_gat) );
AND2XL U_g2046 (.A(G3314_1967_gat), .B(G3344_1970_gat), .Y(G3444_2246_gat) );
AND2XL U_g2047 (.A(G3874_1968_gat), .B(G3989_1969_gat), .Y(G4051_2247_gat) );
BUFX20 U_g2048 (.A(G3874_1968_gat), .Y(G6958_2248_gat) );
BUFX20 U_g2049 (.A(G3874_1968_gat), .Y(G7016_2249_gat) );
AND4XL U_g2050 (.A(G3295_1965_gat), .B(G3335_1113_gat), .C(G3283_1964_gat), .D(G3314_1967_gat), .Y(G3436_2250_gat) );
AND3XL U_g2051 (.A(G3295_1965_gat), .B(G3314_1967_gat), .C(G3335_1113_gat), .Y(G3442_2251_gat) );
AND3XL U_g2052 (.A(G3295_1965_gat), .B(G3335_1113_gat), .C(G3314_1967_gat), .Y(G3439_2252_gat) );
AND2XL U_g2053 (.A(G3335_1113_gat), .B(G3314_1967_gat), .Y(G3443_2253_gat) );
AND2XL U_g2054 (.A(G3335_1113_gat), .B(G3314_1967_gat), .Y(G3445_2254_gat) );
AND3XL U_g2055 (.A(G3856_1966_gat), .B(G3891_1114_gat), .C(G3874_1968_gat), .Y(G4012_2255_gat) );
AND4XL U_g2056 (.A(G3856_1966_gat), .B(G3891_1114_gat), .C(G3845_1963_gat), .D(G3874_1968_gat), .Y(G4009_2256_gat) );
AND3XL U_g2057 (.A(G3856_1966_gat), .B(G3891_1114_gat), .C(G3874_1968_gat), .Y(G4015_2257_gat) );
AND2XL U_g2058 (.A(G3891_1114_gat), .B(G3874_1968_gat), .Y(G4016_2258_gat) );
BUFX20 U_g2059 (.A(G3989_1969_gat), .Y(G7006_2259_gat) );
BUFX20 U_g2060 (.A(G3989_1969_gat), .Y(G6948_2260_gat) );
INVXL U_g2061 (.A(G3344_1970_gat), .Y(G3350_2261_gat) );
BUFX20 U_g2062 (.A(G3899_1971_gat), .Y(G7182_2262_gat) );
BUFX20 U_g2063 (.A(G3899_1971_gat), .Y(G7094_2263_gat) );
AND5XL U_g2064 (.A(G3899_1971_gat), .B(G3911_1974_gat), .C(G3932_1975_gat), .D(G3957_1977_gat), .E(G3997_1980_gat), .Y(G4020_2264_gat) );
AND5XL U_g2065 (.A(G3399_1978_gat), .B(G3353_1972_gat), .C(G3381_1976_gat), .D(G3417_1979_gat), .E(G3365_1973_gat), .Y(G3446_2265_gat) );
BUFX20 U_g2066 (.A(G3353_1972_gat), .Y(G4804_2266_gat) );
AND2XL U_g2067 (.A(G3376_1119_gat), .B(G3353_1972_gat), .Y(G3449_2267_gat) );
AND2XL U_g2068 (.A(G3926_1120_gat), .B(G3899_1971_gat), .Y(G4024_2268_gat) );
BUFX20 U_g2069 (.A(G3365_1973_gat), .Y(G4812_2269_gat) );
BUFX20 U_g2070 (.A(G3911_1974_gat), .Y(G7124_2270_gat) );
AND4XL U_g2071 (.A(G3957_1977_gat), .B(G3911_1974_gat), .C(G3932_1975_gat), .D(G3997_1980_gat), .Y(G4038_2271_gat) );
BUFX20 U_g2072 (.A(G3911_1974_gat), .Y(G7114_2272_gat) );
AND2XL U_g2073 (.A(G3393_1121_gat), .B(G3365_1973_gat), .Y(G3456_2273_gat) );
AND3XL U_g2074 (.A(G3393_1121_gat), .B(G3353_1972_gat), .C(G3365_1973_gat), .Y(G3450_2274_gat) );
AND2XL U_g2075 (.A(G3949_1122_gat), .B(G3911_1974_gat), .Y(G4039_2275_gat) );
AND2XL U_g2076 (.A(G3949_1122_gat), .B(G3911_1974_gat), .Y(G4035_2276_gat) );
AND3XL U_g2077 (.A(G3949_1122_gat), .B(G3899_1971_gat), .C(G3911_1974_gat), .Y(G4025_2277_gat) );
BUFX20 U_g2078 (.A(G3932_1975_gat), .Y(G7192_2278_gat) );
BUFX20 U_g2079 (.A(G3932_1975_gat), .Y(G7104_2279_gat) );
AND3XL U_g2080 (.A(G3957_1977_gat), .B(G3932_1975_gat), .C(G3997_1980_gat), .Y(G4044_2280_gat) );
BUFX20 U_g2081 (.A(G3381_1976_gat), .Y(G4820_2281_gat) );
AND3XL U_g2082 (.A(G3365_1973_gat), .B(G3410_1123_gat), .C(G3381_1976_gat), .Y(G3457_2282_gat) );
AND4XL U_g2083 (.A(G3365_1973_gat), .B(G3410_1123_gat), .C(G3353_1972_gat), .D(G3381_1976_gat), .Y(G3451_2283_gat) );
AND2XL U_g2084 (.A(G3381_1976_gat), .B(G3410_1123_gat), .Y(G3460_2284_gat) );
AND3XL U_g2085 (.A(G3911_1974_gat), .B(G3971_1124_gat), .C(G3932_1975_gat), .Y(G4040_2285_gat) );
AND3XL U_g2086 (.A(G3911_1974_gat), .B(G3971_1124_gat), .C(G3932_1975_gat), .Y(G4036_2286_gat) );
AND4XL U_g2087 (.A(G3911_1974_gat), .B(G3971_1124_gat), .C(G3899_1971_gat), .D(G3932_1975_gat), .Y(G4026_2287_gat) );
AND2XL U_g2088 (.A(G3971_1124_gat), .B(G3932_1975_gat), .Y(G4045_2288_gat) );
AND2XL U_g2089 (.A(G3971_1124_gat), .B(G3932_1975_gat), .Y(G4042_2289_gat) );
BUFX20 U_g2090 (.A(G3957_1977_gat), .Y(G7084_2290_gat) );
BUFX20 U_g2091 (.A(G3957_1977_gat), .Y(G7172_2291_gat) );
AND2XL U_g2092 (.A(G3957_1977_gat), .B(G3997_1980_gat), .Y(G4052_2292_gat) );
BUFX20 U_g2093 (.A(G3399_1978_gat), .Y(G4828_2293_gat) );
AND4XL U_g2094 (.A(G3365_1973_gat), .B(G3425_1125_gat), .C(G3381_1976_gat), .D(G3399_1978_gat), .Y(G3458_2294_gat) );
AND5XL U_g2095 (.A(G3365_1973_gat), .B(G3425_1125_gat), .C(G3353_1972_gat), .D(G3381_1976_gat), .E(G3399_1978_gat), .Y(G3452_2295_gat) );
AND2XL U_g2096 (.A(G3425_1125_gat), .B(G3399_1978_gat), .Y(G3463_2296_gat) );
AND3XL U_g2097 (.A(G3425_1125_gat), .B(G3381_1976_gat), .C(G3399_1978_gat), .Y(G3461_2297_gat) );
AND4XL U_g2098 (.A(G3911_1974_gat), .B(G3979_1126_gat), .C(G3932_1975_gat), .D(G3957_1977_gat), .Y(G4037_2298_gat) );
AND5XL U_g2099 (.A(G3911_1974_gat), .B(G3979_1126_gat), .C(G3899_1971_gat), .D(G3932_1975_gat), .E(G3957_1977_gat), .Y(G4027_2299_gat) );
AND4XL U_g2100 (.A(G3911_1974_gat), .B(G3979_1126_gat), .C(G3932_1975_gat), .D(G3957_1977_gat), .Y(G4041_2300_gat) );
AND3XL U_g2101 (.A(G3979_1126_gat), .B(G3932_1975_gat), .C(G3957_1977_gat), .Y(G4043_2301_gat) );
AND2XL U_g2102 (.A(G3979_1126_gat), .B(G3957_1977_gat), .Y(G4047_2302_gat) );
AND3XL U_g2103 (.A(G3979_1126_gat), .B(G3932_1975_gat), .C(G3957_1977_gat), .Y(G4046_2303_gat) );
BUFX20 U_g2104 (.A(G3417_1979_gat), .Y(G4796_2304_gat) );
BUFX20 U_g2105 (.A(G3997_1980_gat), .Y(G7162_2305_gat) );
BUFX20 U_g2106 (.A(G3997_1980_gat), .Y(G7074_2306_gat) );
AND4XL U_g2107 (.A(G2589_1981_gat), .B(G2600_1984_gat), .C(G2618_1985_gat), .D(G2734_1987_gat), .Y(G2749_2307_gat) );
BUFX20 U_g2108 (.A(G2589_1981_gat), .Y(G6158_2308_gat) );
BUFX20 U_g2109 (.A(G2589_1981_gat), .Y(G6100_2309_gat) );
BUFX20 U_g2110 (.A(G2343_1982_gat), .Y(G5940_2310_gat) );
BUFX20 U_g2111 (.A(G2343_1982_gat), .Y(G5948_2311_gat) );
AND4XL U_g2112 (.A(G2343_1982_gat), .B(G2372_1986_gat), .C(G2400_1988_gat), .D(G2354_1983_gat), .Y(G2487_2312_gat) );
AND2XL U_g2113 (.A(G2366_1130_gat), .B(G2343_1982_gat), .Y(G2492_2313_gat) );
AND2XL U_g2114 (.A(G2612_1131_gat), .B(G2589_1981_gat), .Y(G2754_2314_gat) );
BUFX20 U_g2115 (.A(G2354_1983_gat), .Y(G5964_2315_gat) );
BUFX20 U_g2116 (.A(G2354_1983_gat), .Y(G5956_2316_gat) );
AND3XL U_g2117 (.A(G2354_1983_gat), .B(G2372_1986_gat), .C(G2400_1988_gat), .Y(G2502_2317_gat) );
BUFX20 U_g2118 (.A(G2600_1984_gat), .Y(G6110_2318_gat) );
AND3XL U_g2119 (.A(G2600_1984_gat), .B(G2618_1985_gat), .C(G2734_1987_gat), .Y(G2764_2319_gat) );
BUFX20 U_g2120 (.A(G2600_1984_gat), .Y(G6168_2320_gat) );
AND3XL U_g2121 (.A(G2384_1132_gat), .B(G2343_1982_gat), .C(G2354_1983_gat), .Y(G2493_2321_gat) );
AND2XL U_g2122 (.A(G2384_1132_gat), .B(G2354_1983_gat), .Y(G2500_2322_gat) );
AND2XL U_g2123 (.A(G2384_1132_gat), .B(G2354_1983_gat), .Y(G2503_2323_gat) );
AND2XL U_g2124 (.A(G2629_1133_gat), .B(G2600_1984_gat), .Y(G2765_2324_gat) );
AND3XL U_g2125 (.A(G2629_1133_gat), .B(G2589_1981_gat), .C(G2600_1984_gat), .Y(G2755_2325_gat) );
AND2XL U_g2126 (.A(G2629_1133_gat), .B(G2600_1984_gat), .Y(G2762_2326_gat) );
AND2XL U_g2127 (.A(G2618_1985_gat), .B(G2734_1987_gat), .Y(G2804_2327_gat) );
BUFX20 U_g2128 (.A(G2618_1985_gat), .Y(G6090_2328_gat) );
BUFX20 U_g2129 (.A(G2618_1985_gat), .Y(G6148_2329_gat) );
BUFX20 U_g2130 (.A(G2372_1986_gat), .Y(G5980_2330_gat) );
BUFX20 U_g2131 (.A(G2372_1986_gat), .Y(G5972_2331_gat) );
AND2XL U_g2132 (.A(G2372_1986_gat), .B(G2400_1988_gat), .Y(G2506_2332_gat) );
AND4XL U_g2133 (.A(G2354_1983_gat), .B(G2391_1134_gat), .C(G2343_1982_gat), .D(G2372_1986_gat), .Y(G2494_2333_gat) );
AND3XL U_g2134 (.A(G2354_1983_gat), .B(G2372_1986_gat), .C(G2391_1134_gat), .Y(G2504_2334_gat) );
AND3XL U_g2135 (.A(G2354_1983_gat), .B(G2391_1134_gat), .C(G2372_1986_gat), .Y(G2501_2335_gat) );
AND2XL U_g2136 (.A(G2391_1134_gat), .B(G2372_1986_gat), .Y(G2505_2336_gat) );
AND2XL U_g2137 (.A(G2391_1134_gat), .B(G2372_1986_gat), .Y(G2507_2337_gat) );
AND3XL U_g2138 (.A(G2600_1984_gat), .B(G2635_1135_gat), .C(G2618_1985_gat), .Y(G2763_2338_gat) );
AND4XL U_g2139 (.A(G2600_1984_gat), .B(G2635_1135_gat), .C(G2589_1981_gat), .D(G2618_1985_gat), .Y(G2756_2339_gat) );
AND3XL U_g2140 (.A(G2600_1984_gat), .B(G2635_1135_gat), .C(G2618_1985_gat), .Y(G2766_2340_gat) );
AND2XL U_g2141 (.A(G2635_1135_gat), .B(G2618_1985_gat), .Y(G2767_2341_gat) );
BUFX20 U_g2142 (.A(G2734_1987_gat), .Y(G6138_2342_gat) );
BUFX20 U_g2143 (.A(G2734_1987_gat), .Y(G6080_2343_gat) );
INVXL U_g2144 (.A(G2400_1988_gat), .Y(G2406_2344_gat) );
BUFX20 U_g2145 (.A(G2409_1989_gat), .Y(G4844_2345_gat) );
BUFX20 U_g2146 (.A(G2643_1990_gat), .Y(G6314_2346_gat) );
BUFX20 U_g2147 (.A(G2643_1990_gat), .Y(G6226_2347_gat) );
AND2XL U_g2148 (.A(G2431_1140_gat), .B(G2409_1989_gat), .Y(G2511_2348_gat) );
AND2XL U_g2149 (.A(G2670_1141_gat), .B(G2643_1990_gat), .Y(G2776_2349_gat) );
BUFX20 U_g2150 (.A(G2655_1991_gat), .Y(G6256_2350_gat) );
BUFX20 U_g2151 (.A(G2655_1991_gat), .Y(G6246_2351_gat) );
BUFX20 U_g2152 (.A(G2420_1992_gat), .Y(G4852_2352_gat) );
AND2XL U_g2153 (.A(G2448_1142_gat), .B(G2420_1992_gat), .Y(G2518_2353_gat) );
AND3XL U_g2154 (.A(G2448_1142_gat), .B(G2409_1989_gat), .C(G2420_1992_gat), .Y(G2512_2354_gat) );
AND2XL U_g2155 (.A(G2693_1143_gat), .B(G2655_1991_gat), .Y(G2792_2355_gat) );
AND2XL U_g2156 (.A(G2693_1143_gat), .B(G2655_1991_gat), .Y(G2788_2356_gat) );
AND3XL U_g2157 (.A(G2693_1143_gat), .B(G2643_1990_gat), .C(G2655_1991_gat), .Y(G2777_2357_gat) );
BUFX20 U_g2158 (.A(G2436_1993_gat), .Y(G4860_2358_gat) );
BUFX20 U_g2159 (.A(G2676_1994_gat), .Y(G6324_2359_gat) );
BUFX20 U_g2160 (.A(G2676_1994_gat), .Y(G6236_2360_gat) );
AND3XL U_g2161 (.A(G2420_1992_gat), .B(G2465_1144_gat), .C(G2436_1993_gat), .Y(G2519_2361_gat) );
AND4XL U_g2162 (.A(G2420_1992_gat), .B(G2465_1144_gat), .C(G2409_1989_gat), .D(G2436_1993_gat), .Y(G2513_2362_gat) );
AND2XL U_g2163 (.A(G2436_1993_gat), .B(G2465_1144_gat), .Y(G2523_2363_gat) );
AND3XL U_g2164 (.A(G2655_1991_gat), .B(G2715_1145_gat), .C(G2676_1994_gat), .Y(G2793_2364_gat) );
AND3XL U_g2165 (.A(G2655_1991_gat), .B(G2715_1145_gat), .C(G2676_1994_gat), .Y(G2789_2365_gat) );
AND4XL U_g2166 (.A(G2655_1991_gat), .B(G2715_1145_gat), .C(G2643_1990_gat), .D(G2676_1994_gat), .Y(G2778_2366_gat) );
AND2XL U_g2167 (.A(G2715_1145_gat), .B(G2676_1994_gat), .Y(G2798_2367_gat) );
AND2XL U_g2168 (.A(G2715_1145_gat), .B(G2676_1994_gat), .Y(G2795_2368_gat) );
BUFX20 U_g2169 (.A(G2701_1995_gat), .Y(G6216_2369_gat) );
BUFX20 U_g2170 (.A(G2701_1995_gat), .Y(G6304_2370_gat) );
BUFX20 U_g2171 (.A(G2454_1996_gat), .Y(G4868_2371_gat) );
OR4XL U_g2172 (.A(G3027_2040_gat), .B(G3026_2020_gat), .C(G3025_2005_gat), .D(G2962_867_gat), .Y(G3028_2372_gat) );
OR2XL U_g2173 (.A(G7602_2021_ngat), .B(G7595_1801_ngat), .Y(G7437_2373_gat) );
AND2XL U_g2174 (.A(G3029_2043_gat), .B(G3022_1998_gat), .Y(G3035_2374_gat) );
AND2XL U_g2175 (.A(G1718_2046_gat), .B(G1702_1999_gat), .Y(G1788_2375_gat) );
INVXL U_g2176 (.A(G5566_2000_gat), .Y(G5570_2376_gat) );
INVXL U_g2177 (.A(G5508_2001_gat), .Y(G5512_2377_gat) );
OR4XL U_g2178 (.A(G1707_2029_gat), .B(G1706_2015_gat), .C(G1705_2010_gat), .D(G1553_870_gat), .Y(G1708_2378_gat) );
OR4XL U_g2179 (.A(G1940_2032_gat), .B(G1939_2017_gat), .C(G1938_2006_gat), .D(G1802_871_gat), .Y(G1941_2379_gat) );
INVXL U_g2180 (.A(G5820_2002_gat), .Y(G5824_2380_gat) );
INVXL U_g2181 (.A(G5828_2003_gat), .Y(G5832_2381_gat) );
AND2XL U_g2182 (.A(G1950_2047_gat), .B(G1935_2004_gat), .Y(G1974_2382_gat) );
AND3XL U_g2183 (.A(G1946_2033_ngat), .B(G1945_2019_ngat), .C(G1816_875_ngat), .Y(G5825_2383_gat) );
OR4XL U_g2184 (.A(G1944_2009_gat), .B(G1943_2034_gat), .C(G1942_2018_gat), .D(G1816_875_gat), .Y(G5817_2384_gat) );
INVXL U_g2185 (.A(G5844_2007_gat), .Y(G5848_2385_gat) );
INVXL U_g2186 (.A(G5836_2008_gat), .Y(G5840_2386_gat) );
AND3XL U_g2187 (.A(G1713_2030_ngat), .B(G1712_2014_ngat), .C(G1567_876_ngat), .Y(G5536_2387_gat) );
OR4XL U_g2188 (.A(G1711_2012_gat), .B(G1710_2028_gat), .C(G1709_2016_gat), .D(G1567_876_gat), .Y(G5478_2388_gat) );
INVXL U_g2189 (.A(G5518_2011_gat), .Y(G5522_2389_gat) );
INVXL U_g2190 (.A(G5576_2013_gat), .Y(G5580_2390_gat) );
OR2XL U_g2191 (.A(G1714_2031_gat), .B(G1584_877_gat), .Y(G1715_2391_gat) );
AND2XL U_g2192 (.A(G1949_2036_ngat), .B(G1834_878_ngat), .Y(G5841_2392_gat) );
OR3XL U_g2193 (.A(G1948_2027_gat), .B(G1947_2035_gat), .C(G1834_878_gat), .Y(G5833_2393_gat) );
OR2XL U_g2194 (.A(G7601_1997_ngat), .B(G7598_1809_ngat), .Y(G7436_2394_gat) );
INVXL U_g2195 (.A(G5498_2023_gat), .Y(G5502_2395_gat) );
INVXL U_g2196 (.A(G5556_2024_gat), .Y(G5560_2396_gat) );
INVXL U_g2197 (.A(G5860_2025_gat), .Y(G5864_2397_gat) );
INVXL U_g2198 (.A(G5852_2026_gat), .Y(G5856_2398_gat) );
OR2XL U_g2199 (.A(G5863_1520_ngat), .B(G5860_2025_ngat), .Y(G2003_2399_gat) );
OR2XL U_g2200 (.A(G5855_1161_ngat), .B(G5852_2026_ngat), .Y(G1999_2400_gat) );
INVXL U_g2201 (.A(G5546_2038_gat), .Y(G5550_2401_gat) );
INVXL U_g2202 (.A(G5488_2039_gat), .Y(G5492_2402_gat) );
OR5XL U_g2203 (.A(G3033_2092_gat), .B(G3032_2079_gat), .C(G3031_2061_gat), .D(G3030_2055_gat), .E(G2989_889_gat), .Y(G3034_2403_gat) );
AND3XL U_g2204 (.A(G4602_2041_gat), .B(G4535_2093_gat), .C(G4544_2062_gat), .Y(G4626_2404_gat) );
INVXL U_g2205 (.A(G4602_2041_gat), .Y(G4605_2405_gat) );
INVXL U_g2206 (.A(G4598_2042_gat), .Y(G4601_2406_gat) );
OR5XL U_g2207 (.A(G1725_2081_gat), .B(G1724_2069_gat), .C(G1723_2058_gat), .D(G1722_2049_gat), .E(G1606_892_gat), .Y(G1726_2407_gat) );
INVXL U_g2208 (.A(G5722_2044_gat), .Y(G5726_2408_gat) );
INVXL U_g2209 (.A(G5634_2045_gat), .Y(G5638_2409_gat) );
INVXL U_g2210 (.A(G1718_2046_gat), .Y(G1721_2410_gat) );
OR5XL U_g2211 (.A(G1956_2087_gat), .B(G1955_2073_gat), .C(G1954_2060_gat), .D(G1953_2050_gat), .E(G1866_893_gat), .Y(G1957_2411_gat) );
INVXL U_g2212 (.A(G4724_2048_gat), .Y(G4728_2412_gat) );
AND4XL U_g2213 (.A(G1739_2082_ngat), .B(G1738_2067_ngat), .C(G1737_2056_ngat), .D(G1624_894_ngat), .Y(G5692_2413_gat) );
OR5XL U_g2214 (.A(G1736_2053_gat), .B(G1735_2080_gat), .C(G1734_2068_gat), .D(G1733_2057_gat), .E(G1624_894_gat), .Y(G5604_2414_gat) );
INVXL U_g2215 (.A(G4732_2051_gat), .Y(G4736_2415_gat) );
INVXL U_g2216 (.A(G5664_2052_gat), .Y(G5668_2416_gat) );
INVXL U_g2217 (.A(G5654_2054_gat), .Y(G5658_2417_gat) );
AND3XL U_g2218 (.A(G1744_2085_ngat), .B(G1743_2070_ngat), .C(G1647_899_ngat), .Y(G5672_2418_gat) );
OR4XL U_g2219 (.A(G1742_2065_gat), .B(G1741_2083_gat), .C(G1740_2071_gat), .D(G1647_899_gat), .Y(G5584_2419_gat) );
AND3XL U_g2220 (.A(G4598_2042_gat), .B(G4531_1830_gat), .C(G4540_1822_gat), .Y(G4623_2420_gat) );
INVXL U_g2221 (.A(G5732_2063_gat), .Y(G5736_2421_gat) );
INVXL U_g2222 (.A(G5644_2064_gat), .Y(G5648_2422_gat) );
INVXL U_g2223 (.A(G4740_2066_gat), .Y(G4744_2423_gat) );
OR2XL U_g2224 (.A(G1745_2084_gat), .B(G1669_904_gat), .Y(G1746_2424_gat) );
INVXL U_g2225 (.A(G4748_2075_gat), .Y(G4752_2425_gat) );
INVXL U_g2226 (.A(G5624_2076_gat), .Y(G5628_2426_gat) );
INVXL U_g2227 (.A(G5712_2077_gat), .Y(G5716_2427_gat) );
INVXL U_g2228 (.A(G5702_2090_gat), .Y(G5706_2428_gat) );
INVXL U_g2229 (.A(G5614_2091_gat), .Y(G5618_2429_gat) );
INVXL U_g2230 (.A(G4716_2094_gat), .Y(G4720_2430_gat) );
AND2XL U_g2231 (.A(G1122_2101_gat), .B(G1108_1196_gat), .Y(G1146_2431_gat) );
AND2XL U_g2232 (.A(G920_2100_gat), .B(G902_1199_gat), .Y(G997_2432_gat) );
OR5XL U_g2233 (.A(G928_2126_gat), .B(G927_2112_gat), .C(G926_2163_gat), .D(G925_2103_gat), .E(G802_924_gat), .Y(G929_2433_gat) );
OR5XL U_g2234 (.A(G1128_2132_gat), .B(G1127_2116_gat), .C(G1126_2165_gat), .D(G1125_2104_gat), .E(G1035_925_gat), .Y(G1129_2434_gat) );
OR5XL U_g2235 (.A(G3234_2137_gat), .B(G3233_2119_gat), .C(G3232_2169_gat), .D(G3231_2109_gat), .E(G3183_926_gat), .Y(G3235_2435_gat) );
AND3XL U_g2236 (.A(G3575_2095_gat), .B(G3508_2138_gat), .C(G3517_2120_gat), .Y(G3599_2436_gat) );
INVXL U_g2237 (.A(G3575_2095_gat), .Y(G3578_2437_gat) );
INVXL U_g2238 (.A(G3571_2096_gat), .Y(G3574_2438_gat) );
INVXL U_g2239 (.A(G5152_2098_gat), .Y(G5156_2439_gat) );
INVXL U_g2240 (.A(G5064_2099_gat), .Y(G5068_2440_gat) );
INVXL U_g2241 (.A(G920_2100_gat), .Y(G924_2441_gat) );
INVXL U_g2242 (.A(G4764_2102_gat), .Y(G4768_2442_gat) );
AND4XL U_g2243 (.A(G943_2127_ngat), .B(G942_2110_ngat), .C(G941_2161_ngat), .D(G821_929_ngat), .Y(G5122_2443_gat) );
OR5XL U_g2244 (.A(G940_2107_gat), .B(G939_2125_gat), .C(G938_2111_gat), .D(G937_2162_gat), .E(G821_929_gat), .Y(G5034_2444_gat) );
INVXL U_g2245 (.A(G4772_2105_gat), .Y(G4776_2445_gat) );
INVXL U_g2246 (.A(G5094_2106_gat), .Y(G5098_2446_gat) );
INVXL U_g2247 (.A(G5084_2108_gat), .Y(G5088_2447_gat) );
OR2XL U_g2248 (.A(G949_2129_gat), .B(G868_934_gat), .Y(G950_2448_gat) );
INVXL U_g2249 (.A(G4788_2118_gat), .Y(G4792_2449_gat) );
AND3XL U_g2250 (.A(G3571_2096_gat), .B(G3504_1851_gat), .C(G3513_1848_gat), .Y(G3596_2450_gat) );
INVXL U_g2251 (.A(G5054_2121_gat), .Y(G5058_2451_gat) );
INVXL U_g2252 (.A(G5142_2123_gat), .Y(G5146_2452_gat) );
INVXL U_g2253 (.A(G5132_2135_gat), .Y(G5136_2453_gat) );
INVXL U_g2254 (.A(G5044_2136_gat), .Y(G5048_2454_gat) );
INVXL U_g2255 (.A(G4756_2139_gat), .Y(G4760_2455_gat) );
AND3XL U_g2256 (.A(G4263_2142_gat), .B(G4226_1854_gat), .C(G4235_1855_gat), .Y(G4284_2456_gat) );
AND3XL U_g2257 (.A(G4267_2143_gat), .B(G4230_2140_gat), .C(G4239_2141_gat), .Y(G4287_2457_gat) );
INVXL U_g2258 (.A(G4263_2142_gat), .Y(G4266_2458_gat) );
INVXL U_g2259 (.A(G4267_2143_gat), .Y(G4270_2459_gat) );
AND3XL U_g2260 (.A(G1300_2146_gat), .B(G1263_1857_gat), .C(G1272_1858_gat), .Y(G1321_2460_gat) );
AND3XL U_g2261 (.A(G1304_2147_gat), .B(G1267_2144_gat), .C(G1276_2145_gat), .Y(G1324_2461_gat) );
INVXL U_g2262 (.A(G1300_2146_gat), .Y(G1303_2462_gat) );
INVXL U_g2263 (.A(G1304_2147_gat), .Y(G1307_2463_gat) );
INVXL U_g2264 (.A(G7348_2148_gat), .Y(G7352_2464_gat) );
AND4XL U_g2265 (.A(G4300_2153_gat), .B(G4314_1248_gat), .C(G4291_2173_gat), .D(G4308_2151_gat), .Y(G4363_2465_gat) );
AND4XL U_g2266 (.A(G4291_2173_gat), .B(G4300_2153_gat), .C(G4308_2151_gat), .D(G4352_2149_gat), .Y(G4356_2466_gat) );
INVXL U_g2267 (.A(G6822_2150_gat), .Y(G6826_2467_gat) );
AND3XL U_g2268 (.A(G4312_1256_gat), .B(G4291_2173_gat), .C(G4300_2153_gat), .Y(G4362_2468_gat) );
INVXL U_g2269 (.A(G6819_2152_gat), .Y(G6825_2469_gat) );
AND2XL U_g2270 (.A(G4305_1262_gat), .B(G4291_2173_gat), .Y(G4361_2470_gat) );
INVXL U_g2271 (.A(G7345_2154_gat), .Y(G7351_2471_gat) );
BUFX20 U_g2272 (.A(G3545_2155_gat), .Y(G3583_2472_gat) );
BUFX20 U_g2273 (.A(G3545_2155_gat), .Y(G3579_2473_gat) );
AND2XL U_g2274 (.A(G3099_1268_gat), .B(G3082_2179_gat), .Y(G3139_2474_gat) );
AND5XL U_g2275 (.A(G3082_2179_gat), .B(G3093_2156_gat), .C(G3102_2177_gat), .D(G3110_2175_gat), .E(G3122_2158_gat), .Y(G3136_2475_gat) );
BUFX20 U_g2276 (.A(G4198_2157_gat), .Y(G4251_2476_gat) );
BUFX20 U_g2277 (.A(G4198_2157_gat), .Y(G4247_2477_gat) );
AND5XL U_g2278 (.A(G3093_2156_gat), .B(G3116_1271_gat), .C(G3082_2179_gat), .D(G3102_2177_gat), .E(G3110_2175_gat), .Y(G3142_2478_gat) );
INVXL U_g2279 (.A(G4180_2159_gat), .Y(G4184_2479_gat) );
INVXL U_g2280 (.A(G3527_2160_gat), .Y(G3531_2480_gat) );
AND3XL U_g2281 (.A(G948_2130_ngat), .B(G947_2113_ngat), .C(G845_980_ngat), .Y(G5102_2481_gat) );
OR4XL U_g2282 (.A(G946_2122_gat), .B(G945_2128_gat), .C(G944_2114_gat), .D(G845_980_gat), .Y(G5014_2482_gat) );
INVXL U_g2283 (.A(G5162_2166_gat), .Y(G5166_2483_gat) );
INVXL U_g2284 (.A(G5074_2167_gat), .Y(G5078_2484_gat) );
INVXL U_g2285 (.A(G4780_2168_gat), .Y(G4784_2485_gat) );
AND5XL U_g2286 (.A(G4317_2170_gat), .B(G4327_2186_gat), .C(G4336_2185_gat), .D(G4344_2188_gat), .E(G4355_2207_gat), .Y(G4369_2486_gat) );
BUFX20 U_g2287 (.A(G4221_2171_gat), .Y(G4259_2487_gat) );
BUFX20 U_g2288 (.A(G4221_2171_gat), .Y(G4255_2488_gat) );
BUFX20 U_g2289 (.A(G3568_2172_gat), .Y(G3587_2489_gat) );
BUFX20 U_g2290 (.A(G3568_2172_gat), .Y(G3591_2490_gat) );
INVXL U_g2291 (.A(G3536_2174_gat), .Y(G3540_2491_gat) );
AND4XL U_g2292 (.A(G3093_2156_gat), .B(G3114_1298_gat), .C(G3082_2179_gat), .D(G3102_2177_gat), .Y(G3141_2492_gat) );
INVXL U_g2293 (.A(G4189_2176_gat), .Y(G4193_2493_gat) );
AND3XL U_g2294 (.A(G3107_1305_gat), .B(G3082_2179_gat), .C(G3093_2156_gat), .Y(G3140_2494_gat) );
BUFX20 U_g2295 (.A(G4595_2178_gat), .Y(G4614_2495_gat) );
BUFX20 U_g2296 (.A(G4595_2178_gat), .Y(G4618_2496_gat) );
AND4XL U_g2297 (.A(G3052_2192_gat), .B(G3062_2194_gat), .C(G3071_2195_gat), .D(G3119_2180_gat), .Y(G3123_2497_gat) );
INVXL U_g2298 (.A(G7614_2181_gat), .Y(G7618_2498_gat) );
INVXL U_g2299 (.A(G4586_2182_gat), .Y(G4590_2499_gat) );
INVXL U_g2300 (.A(G4577_2183_gat), .Y(G4581_2500_gat) );
INVXL U_g2301 (.A(G4563_2184_gat), .Y(G4567_2501_gat) );
BUFX20 U_g2302 (.A(G4572_2187_gat), .Y(G4610_2502_gat) );
BUFX20 U_g2303 (.A(G4572_2187_gat), .Y(G4606_2503_gat) );
INVXL U_g2304 (.A(G6809_2190_gat), .Y(G6815_2504_gat) );
OR2XL U_g2305 (.A(G7344_2203_ngat), .B(G7337_1902_ngat), .Y(G6351_2505_gat) );
INVXL U_g2306 (.A(G7611_2193_gat), .Y(G7617_2506_gat) );
INVXL U_g2307 (.A(G7603_2196_gat), .Y(G7609_2507_gat) );
INVXL U_g2308 (.A(G7606_2197_gat), .Y(G7610_2508_gat) );
AND2XL U_g2309 (.A(G3068_1353_gat), .B(G3052_2192_gat), .Y(G3128_2509_gat) );
INVXL U_g2310 (.A(G3550_2199_gat), .Y(G3554_2510_gat) );
OR2XL U_g2311 (.A(G4979_2200_ngat), .B(G4978_1926_ngat), .Y(G4980_2511_gat) );
OR2XL U_g2312 (.A(G4938_2202_ngat), .B(G4937_1929_ngat), .Y(G4939_2512_gat) );
AND4XL U_g2313 (.A(G3062_2194_gat), .B(G3079_1370_gat), .C(G3052_2192_gat), .D(G3071_2195_gat), .Y(G3130_2513_gat) );
OR2XL U_g2314 (.A(G7343_2191_ngat), .B(G7340_1931_ngat), .Y(G6350_2514_gat) );
INVXL U_g2315 (.A(G6812_2204_gat), .Y(G6816_2515_gat) );
AND3XL U_g2316 (.A(G3076_1379_gat), .B(G3052_2192_gat), .C(G3062_2194_gat), .Y(G3129_2516_gat) );
INVXL U_g2317 (.A(G3559_2205_gat), .Y(G3563_2517_gat) );
AND4XL U_g2318 (.A(G4327_2186_gat), .B(G4348_1385_gat), .C(G4317_2170_gat), .D(G4336_2185_gat), .Y(G4374_2518_gat) );
AND3XL U_g2319 (.A(G4341_1392_gat), .B(G4317_2170_gat), .C(G4327_2186_gat), .Y(G4373_2519_gat) );
AND2XL U_g2320 (.A(G4333_1397_gat), .B(G4317_2170_gat), .Y(G4372_2520_gat) );
AND5XL U_g2321 (.A(G4327_2186_gat), .B(G4349_1400_gat), .C(G4317_2170_gat), .D(G4336_2185_gat), .E(G4344_2188_gat), .Y(G4375_2521_gat) );
AND4XL U_g2322 (.A(G2420_1992_gat), .B(G2481_1721_gat), .C(G2436_1993_gat), .D(G2454_1996_gat), .Y(G2520_2522_gat) );
AND5XL U_g2323 (.A(G2420_1992_gat), .B(G2481_1721_gat), .C(G2409_1989_gat), .D(G2436_1993_gat), .E(G2454_1996_gat), .Y(G2514_2523_gat) );
AND2XL U_g2324 (.A(G2481_1721_gat), .B(G2454_1996_gat), .Y(G2527_2524_gat) );
AND3XL U_g2325 (.A(G2481_1721_gat), .B(G2436_1993_gat), .C(G2454_1996_gat), .Y(G2524_2525_gat) );
AND4XL U_g2326 (.A(G2655_1991_gat), .B(G2724_1722_gat), .C(G2676_1994_gat), .D(G2701_1995_gat), .Y(G2790_2526_gat) );
AND5XL U_g2327 (.A(G2655_1991_gat), .B(G2724_1722_gat), .C(G2643_1990_gat), .D(G2676_1994_gat), .E(G2701_1995_gat), .Y(G2779_2527_gat) );
AND4XL U_g2328 (.A(G2655_1991_gat), .B(G2724_1722_gat), .C(G2676_1994_gat), .D(G2701_1995_gat), .Y(G2794_2528_gat) );
AND3XL U_g2329 (.A(G2724_1722_gat), .B(G2676_1994_gat), .C(G2701_1995_gat), .Y(G2796_2529_gat) );
AND2XL U_g2330 (.A(G2724_1722_gat), .B(G2701_1995_gat), .Y(G2800_2530_gat) );
AND3XL U_g2331 (.A(G2724_1722_gat), .B(G2676_1994_gat), .C(G2701_1995_gat), .Y(G2799_2531_gat) );
OR2XL U_g2332 (.A(G2471_2209_ngat), .B(G2470_1945_ngat), .Y(G2472_2532_gat) );
OR2XL U_g2333 (.A(G2741_2210_ngat), .B(G2740_1947_ngat), .Y(G2742_2533_gat) );
AND3XL U_g2334 (.A(G1292_2213_gat), .B(G1240_1950_gat), .C(G1249_1952_gat), .Y(G1315_2534_gat) );
AND3XL U_g2335 (.A(G1296_2212_gat), .B(G1244_2211_gat), .C(G1253_2214_gat), .Y(G1318_2535_gat) );
INVXL U_g2336 (.A(G1296_2212_gat), .Y(G1299_2536_gat) );
INVXL U_g2337 (.A(G1292_2213_gat), .Y(G1295_2537_gat) );
OR2XL U_g2338 (.A(G7360_2216_ngat), .B(G7353_1954_ngat), .Y(G6341_2538_gat) );
OR2XL U_g2339 (.A(G7359_2215_ngat), .B(G7356_1955_ngat), .Y(G6340_2539_gat) );
OR2XL U_g2340 (.A(G5365_2218_ngat), .B(G5362_1956_ngat), .Y(G5367_2540_gat) );
OR2XL U_g2341 (.A(G5366_2217_ngat), .B(G5359_1957_ngat), .Y(G5368_2541_gat) );
AND3XL U_g2342 (.A(G1288_2219_gat), .B(G1221_2222_gat), .C(G1230_2221_gat), .Y(G1312_2542_gat) );
INVXL U_g2343 (.A(G1288_2219_gat), .Y(G1291_2543_gat) );
INVXL U_g2344 (.A(G1284_2220_gat), .Y(G1287_2544_gat) );
AND3XL U_g2345 (.A(G1284_2220_gat), .B(G1217_1960_gat), .C(G1226_1959_gat), .Y(G1309_2545_gat) );
AND2XL U_g2346 (.A(G3235_2435_gat), .B(G3216_1462_gat), .Y(G3258_2546_gat) );
AND2XL U_g2347 (.A(G2472_2532_gat), .B(G4526_205_gat), .Y(G2531_2547_gat) );
AND3XL U_g2348 (.A(G2454_1996_gat), .B(G2472_2532_gat), .C(G4526_205_gat), .Y(G2529_2548_gat) );
AND4XL U_g2349 (.A(G2454_1996_gat), .B(G2436_1993_gat), .C(G2472_2532_gat), .D(G4526_205_gat), .Y(G2526_2549_gat) );
AND5XL U_g2350 (.A(G2420_1992_gat), .B(G2454_1996_gat), .C(G2436_1993_gat), .D(G2472_2532_gat), .E(G4526_205_gat), .Y(G2522_2550_gat) );
OR4XL U_g2351 (.A(G3436_2250_gat), .B(G3435_2238_gat), .C(G3434_2230_gat), .D(G3292_1107_gat), .Y(G3437_2551_gat) );
OR4XL U_g2352 (.A(G4009_2256_gat), .B(G4008_2242_gat), .C(G4007_2231_gat), .D(G3853_1108_gat), .Y(G4010_2552_gat) );
AND2XL U_g2353 (.A(G4020_2264_gat), .B(G4004_2224_gat), .Y(G4089_2553_gat) );
INVXL U_g2354 (.A(G7026_2225_gat), .Y(G7030_2554_gat) );
INVXL U_g2355 (.A(G6968_2226_gat), .Y(G6972_2555_gat) );
INVXL U_g2356 (.A(G6642_2227_gat), .Y(G6646_2556_gat) );
INVXL U_g2357 (.A(G6650_2228_gat), .Y(G6654_2557_gat) );
AND2XL U_g2358 (.A(G3446_2265_gat), .B(G3431_2229_gat), .Y(G3466_2558_gat) );
AND3XL U_g2359 (.A(G3442_2251_ngat), .B(G3441_2240_ngat), .C(G3308_1109_ngat), .Y(G6647_2559_gat) );
OR4XL U_g2360 (.A(G3440_2234_gat), .B(G3439_2252_gat), .C(G3438_2239_gat), .D(G3308_1109_gat), .Y(G6639_2560_gat) );
AND3XL U_g2361 (.A(G4015_2257_ngat), .B(G4014_2241_ngat), .C(G3868_1110_ngat), .Y(G6996_2561_gat) );
OR4XL U_g2362 (.A(G4013_2236_gat), .B(G4012_2255_gat), .C(G4011_2243_gat), .D(G3868_1110_gat), .Y(G6938_2562_gat) );
INVXL U_g2363 (.A(G6666_2232_gat), .Y(G6670_2563_gat) );
INVXL U_g2364 (.A(G6658_2233_gat), .Y(G6662_2564_gat) );
INVXL U_g2365 (.A(G6978_2235_gat), .Y(G6982_2565_gat) );
INVXL U_g2366 (.A(G7036_2237_gat), .Y(G7040_2566_gat) );
AND2XL U_g2367 (.A(G3445_2254_ngat), .B(G3327_1111_ngat), .Y(G6663_2567_gat) );
OR3XL U_g2368 (.A(G3444_2246_gat), .B(G3443_2253_gat), .C(G3327_1111_gat), .Y(G6655_2568_gat) );
OR2XL U_g2369 (.A(G4016_2258_gat), .B(G3885_1112_gat), .Y(G4017_2569_gat) );
INVXL U_g2370 (.A(G6682_2244_gat), .Y(G6686_2570_gat) );
INVXL U_g2371 (.A(G6674_2245_gat), .Y(G6678_2571_gat) );
INVXL U_g2372 (.A(G6958_2248_gat), .Y(G6962_2572_gat) );
INVXL U_g2373 (.A(G7016_2249_gat), .Y(G7020_2573_gat) );
OR2XL U_g2374 (.A(G6685_1768_ngat), .B(G6682_2244_ngat), .Y(G3487_2574_gat) );
INVXL U_g2375 (.A(G7006_2259_gat), .Y(G7010_2575_gat) );
INVXL U_g2376 (.A(G6948_2260_gat), .Y(G6952_2576_gat) );
OR2XL U_g2377 (.A(G6677_1474_ngat), .B(G6674_2245_ngat), .Y(G3483_2577_gat) );
OR5XL U_g2378 (.A(G3452_2295_gat), .B(G3451_2283_gat), .C(G3450_2274_gat), .D(G3449_2267_gat), .E(G3362_1117_gat), .Y(G3453_2578_gat) );
OR5XL U_g2379 (.A(G4027_2299_gat), .B(G4026_2287_gat), .C(G4025_2277_gat), .D(G4024_2268_gat), .E(G3908_1118_gat), .Y(G4028_2579_gat) );
INVXL U_g2380 (.A(G7182_2262_gat), .Y(G7186_2580_gat) );
INVXL U_g2381 (.A(G7094_2263_gat), .Y(G7098_2581_gat) );
INVXL U_g2382 (.A(G4020_2264_gat), .Y(G4023_2582_gat) );
INVXL U_g2383 (.A(G4804_2266_gat), .Y(G4808_2583_gat) );
AND4XL U_g2384 (.A(G4041_2300_ngat), .B(G4040_2285_ngat), .C(G4039_2275_ngat), .D(G3926_1120_ngat), .Y(G7152_2584_gat) );
OR5XL U_g2385 (.A(G4038_2271_gat), .B(G4037_2298_gat), .C(G4036_2286_gat), .D(G4035_2276_gat), .E(G3926_1120_gat), .Y(G7064_2585_gat) );
INVXL U_g2386 (.A(G4812_2269_gat), .Y(G4816_2586_gat) );
INVXL U_g2387 (.A(G7124_2270_gat), .Y(G7128_2587_gat) );
INVXL U_g2388 (.A(G7114_2272_gat), .Y(G7118_2588_gat) );
AND3XL U_g2389 (.A(G4046_2303_ngat), .B(G4045_2288_ngat), .C(G3949_1122_ngat), .Y(G7132_2589_gat) );
OR4XL U_g2390 (.A(G4044_2280_gat), .B(G4043_2301_gat), .C(G4042_2289_gat), .D(G3949_1122_gat), .Y(G7044_2590_gat) );
INVXL U_g2391 (.A(G7192_2278_gat), .Y(G7196_2591_gat) );
INVXL U_g2392 (.A(G7104_2279_gat), .Y(G7108_2592_gat) );
INVXL U_g2393 (.A(G4820_2281_gat), .Y(G4824_2593_gat) );
OR2XL U_g2394 (.A(G4047_2302_gat), .B(G3971_1124_gat), .Y(G4048_2594_gat) );
INVXL U_g2395 (.A(G7084_2290_gat), .Y(G7088_2595_gat) );
INVXL U_g2396 (.A(G7172_2291_gat), .Y(G7176_2596_gat) );
INVXL U_g2397 (.A(G4828_2293_gat), .Y(G4832_2597_gat) );
INVXL U_g2398 (.A(G4796_2304_gat), .Y(G4800_2598_gat) );
INVXL U_g2399 (.A(G7162_2305_gat), .Y(G7166_2599_gat) );
INVXL U_g2400 (.A(G7074_2306_gat), .Y(G7078_2600_gat) );
OR4XL U_g2401 (.A(G2494_2333_gat), .B(G2493_2321_gat), .C(G2492_2313_gat), .D(G2351_1128_gat), .Y(G2495_2601_gat) );
OR4XL U_g2402 (.A(G2756_2339_gat), .B(G2755_2325_gat), .C(G2754_2314_gat), .D(G2597_1129_gat), .Y(G2757_2602_gat) );
INVXL U_g2403 (.A(G2749_2307_gat), .Y(G2753_2603_gat) );
INVXL U_g2404 (.A(G6158_2308_gat), .Y(G6162_2604_gat) );
INVXL U_g2405 (.A(G6100_2309_gat), .Y(G6104_2605_gat) );
INVXL U_g2406 (.A(G5940_2310_gat), .Y(G5944_2606_gat) );
INVXL U_g2407 (.A(G5948_2311_gat), .Y(G5952_2607_gat) );
INVXL U_g2408 (.A(G2487_2312_gat), .Y(G2491_2608_gat) );
AND3XL U_g2409 (.A(G2504_2334_ngat), .B(G2503_2323_ngat), .C(G2366_1130_ngat), .Y(G5945_2609_gat) );
OR4XL U_g2410 (.A(G2502_2317_gat), .B(G2501_2335_gat), .C(G2500_2322_gat), .D(G2366_1130_gat), .Y(G5937_2610_gat) );
AND3XL U_g2411 (.A(G2766_2340_ngat), .B(G2765_2324_ngat), .C(G2612_1131_ngat), .Y(G6128_2611_gat) );
OR4XL U_g2412 (.A(G2764_2319_gat), .B(G2763_2338_gat), .C(G2762_2326_gat), .D(G2612_1131_gat), .Y(G6070_2612_gat) );
INVXL U_g2413 (.A(G5964_2315_gat), .Y(G5968_2613_gat) );
INVXL U_g2414 (.A(G5956_2316_gat), .Y(G5960_2614_gat) );
INVXL U_g2415 (.A(G6110_2318_gat), .Y(G6114_2615_gat) );
INVXL U_g2416 (.A(G6168_2320_gat), .Y(G6172_2616_gat) );
AND2XL U_g2417 (.A(G2507_2337_ngat), .B(G2384_1132_ngat), .Y(G5961_2617_gat) );
OR3XL U_g2418 (.A(G2506_2332_gat), .B(G2505_2336_gat), .C(G2384_1132_gat), .Y(G5953_2618_gat) );
OR2XL U_g2419 (.A(G2767_2341_gat), .B(G2629_1133_gat), .Y(G2768_2619_gat) );
INVXL U_g2420 (.A(G6090_2328_gat), .Y(G6094_2620_gat) );
INVXL U_g2421 (.A(G6148_2329_gat), .Y(G6152_2621_gat) );
INVXL U_g2422 (.A(G5980_2330_gat), .Y(G5984_2622_gat) );
INVXL U_g2423 (.A(G5972_2331_gat), .Y(G5976_2623_gat) );
OR2XL U_g2424 (.A(G5983_1789_ngat), .B(G5980_2330_ngat), .Y(G2559_2624_gat) );
INVXL U_g2425 (.A(G6138_2342_gat), .Y(G6142_2625_gat) );
INVXL U_g2426 (.A(G6080_2343_gat), .Y(G6084_2626_gat) );
OR2XL U_g2427 (.A(G5975_1498_ngat), .B(G5972_2331_ngat), .Y(G2555_2627_gat) );
OR5XL U_g2428 (.A(G2514_2523_gat), .B(G2513_2362_gat), .C(G2512_2354_gat), .D(G2511_2348_gat), .E(G2417_1138_gat), .Y(G2515_2628_gat) );
OR5XL U_g2429 (.A(G2779_2527_gat), .B(G2778_2366_gat), .C(G2777_2357_gat), .D(G2776_2349_gat), .E(G2652_1139_gat), .Y(G2780_2629_gat) );
AND5XL U_g2430 (.A(G2454_1996_gat), .B(G2409_1989_gat), .C(G2436_1993_gat), .D(G2472_2532_gat), .E(G2420_1992_gat), .Y(G2508_2630_gat) );
INVXL U_g2431 (.A(G4844_2345_gat), .Y(G4848_2631_gat) );
INVXL U_g2432 (.A(G6314_2346_gat), .Y(G6318_2632_gat) );
INVXL U_g2433 (.A(G6226_2347_gat), .Y(G6230_2633_gat) );
AND5XL U_g2434 (.A(G2643_1990_gat), .B(G2655_1991_gat), .C(G2676_1994_gat), .D(G2701_1995_gat), .E(G2742_2533_gat), .Y(G2771_2634_gat) );
AND4XL U_g2435 (.A(G2794_2528_ngat), .B(G2793_2364_ngat), .C(G2792_2355_ngat), .D(G2670_1141_ngat), .Y(G6284_2635_gat) );
INVXL U_g2436 (.A(G6256_2350_gat), .Y(G6260_2636_gat) );
AND4XL U_g2437 (.A(G2701_1995_gat), .B(G2655_1991_gat), .C(G2676_1994_gat), .D(G2742_2533_gat), .Y(G2791_2637_gat) );
INVXL U_g2438 (.A(G6246_2351_gat), .Y(G6250_2638_gat) );
INVXL U_g2439 (.A(G4852_2352_gat), .Y(G4856_2639_gat) );
AND3XL U_g2440 (.A(G2799_2531_ngat), .B(G2798_2367_ngat), .C(G2693_1143_ngat), .Y(G6264_2640_gat) );
INVXL U_g2441 (.A(G4860_2358_gat), .Y(G4864_2641_gat) );
INVXL U_g2442 (.A(G6324_2359_gat), .Y(G6328_2642_gat) );
INVXL U_g2443 (.A(G6236_2360_gat), .Y(G6240_2643_gat) );
AND3XL U_g2444 (.A(G2701_1995_gat), .B(G2676_1994_gat), .C(G2742_2533_gat), .Y(G2797_2644_gat) );
OR2XL U_g2445 (.A(G2800_2530_gat), .B(G2715_1145_gat), .Y(G2801_2645_gat) );
INVXL U_g2446 (.A(G6216_2369_gat), .Y(G6220_2646_gat) );
INVXL U_g2447 (.A(G6304_2370_gat), .Y(G6308_2647_gat) );
AND2XL U_g2448 (.A(G2701_1995_gat), .B(G2742_2533_gat), .Y(G2807_2648_gat) );
INVXL U_g2449 (.A(G4868_2371_gat), .Y(G4872_2649_gat) );
OR2XL U_g2450 (.A(G7437_2373_ngat), .B(G7436_2394_ngat), .Y(G7438_2650_gat) );
AND2XL U_g2451 (.A(G3034_2403_gat), .B(G3022_1998_gat), .Y(G3045_2651_gat) );
AND2XL U_g2452 (.A(G1726_2407_gat), .B(G1702_1999_gat), .Y(G1789_2652_gat) );
OR2XL U_g2453 (.A(G5824_2380_ngat), .B(G5817_2384_ngat), .Y(G1986_2653_gat) );
OR2XL U_g2454 (.A(G5832_2381_ngat), .B(G5825_2383_ngat), .Y(G1989_2654_gat) );
AND2XL U_g2455 (.A(G1935_2004_gat), .B(G1957_2411_gat), .Y(G1981_2655_gat) );
INVXL U_g2456 (.A(G5825_2383_gat), .Y(G5831_2656_gat) );
INVXL U_g2457 (.A(G5817_2384_gat), .Y(G5823_2657_gat) );
OR2XL U_g2458 (.A(G5848_2385_ngat), .B(G5841_2392_ngat), .Y(G1996_2658_gat) );
OR2XL U_g2459 (.A(G5840_2386_ngat), .B(G5833_2393_ngat), .Y(G1993_2659_gat) );
INVXL U_g2460 (.A(G5536_2387_gat), .Y(G5540_2660_gat) );
INVXL U_g2461 (.A(G5478_2388_gat), .Y(G5482_2661_gat) );
INVXL U_g2462 (.A(G1715_2391_gat), .Y(G5526_2662_gat) );
INVXL U_g2463 (.A(G5841_2392_gat), .Y(G5847_2663_gat) );
INVXL U_g2464 (.A(G5833_2393_gat), .Y(G5839_2664_gat) );
OR2XL U_g2465 (.A(G1749_2022_gat), .B(G1715_2391_gat), .Y(G5468_2665_gat) );
OR2XL U_g2466 (.A(G5864_2397_ngat), .B(G5857_1159_ngat), .Y(G2004_2666_gat) );
OR2XL U_g2467 (.A(G5856_2398_ngat), .B(G5849_884_ngat), .Y(G2000_2667_gat) );
INVXL U_g2468 (.A(G1726_2407_gat), .Y(G1730_2668_gat) );
INVXL U_g2469 (.A(G5692_2413_gat), .Y(G5696_2669_gat) );
INVXL U_g2470 (.A(G5604_2414_gat), .Y(G5608_2670_gat) );
INVXL U_g2471 (.A(G5672_2418_gat), .Y(G5676_2671_gat) );
INVXL U_g2472 (.A(G5584_2419_gat), .Y(G5588_2672_gat) );
AND3XL U_g2473 (.A(G4601_2406_gat), .B(G4540_1822_gat), .C(G4535_2093_gat), .Y(G4622_2673_gat) );
INVXL U_g2474 (.A(G1746_2424_gat), .Y(G5682_2674_gat) );
OR2XL U_g2475 (.A(G1750_2078_gat), .B(G1746_2424_gat), .Y(G5594_2675_gat) );
OR2XL U_g2476 (.A(G5675_1541_ngat), .B(G5672_2418_ngat), .Y(G5677_2676_gat) );
OR2XL U_g2477 (.A(G5587_1183_ngat), .B(G5584_2419_ngat), .Y(G5589_2677_gat) );
AND3XL U_g2478 (.A(G4605_2405_gat), .B(G4544_2062_gat), .C(G4531_1830_gat), .Y(G4625_2678_gat) );
OR2XL U_g2479 (.A(G4987_1549_ngat), .B(G4980_2511_ngat), .Y(G4989_2679_gat) );
OR2XL U_g2480 (.A(G4946_1837_ngat), .B(G4939_2512_ngat), .Y(G4948_2680_gat) );
AND2XL U_g2481 (.A(G1108_1196_gat), .B(G1129_2434_gat), .Y(G1151_2681_gat) );
AND2XL U_g2482 (.A(G929_2433_gat), .B(G902_1199_gat), .Y(G1002_2682_gat) );
INVXL U_g2483 (.A(G929_2433_gat), .Y(G933_2683_gat) );
INVXL U_g2484 (.A(G3235_2435_gat), .Y(G3238_2684_gat) );
INVXL U_g2485 (.A(G5122_2443_gat), .Y(G5126_2685_gat) );
INVXL U_g2486 (.A(G5034_2444_gat), .Y(G5038_2686_gat) );
INVXL U_g2487 (.A(G950_2448_gat), .Y(G5112_2687_gat) );
AND3XL U_g2488 (.A(G3574_2438_gat), .B(G3513_1848_gat), .C(G3508_2138_gat), .Y(G3595_2688_gat) );
OR2XL U_g2489 (.A(G956_2124_gat), .B(G950_2448_gat), .Y(G5024_2689_gat) );
OR2XL U_g2490 (.A(G5105_1569_ngat), .B(G5102_2481_ngat), .Y(G5107_2690_gat) );
OR2XL U_g2491 (.A(G5017_1219_ngat), .B(G5014_2482_ngat), .Y(G5019_2691_gat) );
AND3XL U_g2492 (.A(G3578_2437_gat), .B(G3517_2120_gat), .C(G3504_1851_gat), .Y(G3598_2692_gat) );
AND3XL U_g2493 (.A(G4270_2459_gat), .B(G4239_2141_gat), .C(G4226_1854_gat), .Y(G4286_2693_gat) );
AND3XL U_g2494 (.A(G4266_2458_gat), .B(G4235_1855_gat), .C(G4230_2140_gat), .Y(G4283_2694_gat) );
AND3XL U_g2495 (.A(G1307_2463_gat), .B(G1276_2145_gat), .C(G1263_1857_gat), .Y(G1323_2695_gat) );
AND3XL U_g2496 (.A(G1303_2462_gat), .B(G1272_1858_gat), .C(G1267_2144_gat), .Y(G1320_2696_gat) );
OR2XL U_g2497 (.A(G7351_2471_ngat), .B(G7348_2148_ngat), .Y(G6360_2697_gat) );
AND2XL U_g2498 (.A(G4369_2486_gat), .B(G4356_2466_gat), .Y(G4386_2698_gat) );
INVXL U_g2499 (.A(G4356_2466_gat), .Y(G4360_2699_gat) );
OR2XL U_g2500 (.A(G6825_2469_ngat), .B(G6822_2150_ngat), .Y(G6827_2700_gat) );
OR2XL U_g2501 (.A(G6826_2467_ngat), .B(G6819_2152_ngat), .Y(G6828_2701_gat) );
OR2XL U_g2502 (.A(G7352_2464_ngat), .B(G7345_2154_ngat), .Y(G6361_2702_gat) );
AND3XL U_g2503 (.A(G3583_2472_gat), .B(G3531_2480_gat), .C(G3540_2491_gat), .Y(G3605_2703_gat) );
INVXL U_g2504 (.A(G3583_2472_gat), .Y(G3586_2704_gat) );
INVXL U_g2505 (.A(G3579_2473_gat), .Y(G3582_2705_gat) );
AND2XL U_g2506 (.A(G3136_2475_gat), .B(G3123_2497_gat), .Y(G3156_2706_gat) );
AND3XL U_g2507 (.A(G4251_2476_gat), .B(G4184_2479_gat), .C(G4193_2493_gat), .Y(G4275_2707_gat) );
INVXL U_g2508 (.A(G4251_2476_gat), .Y(G4254_2708_gat) );
INVXL U_g2509 (.A(G4247_2477_gat), .Y(G4250_2709_gat) );
AND3XL U_g2510 (.A(G4247_2477_gat), .B(G4180_2159_gat), .C(G4189_2176_gat), .Y(G4272_2710_gat) );
AND3XL U_g2511 (.A(G3579_2473_gat), .B(G3527_2160_gat), .C(G3536_2174_gat), .Y(G3602_2711_gat) );
INVXL U_g2512 (.A(G5102_2481_gat), .Y(G5106_2712_gat) );
INVXL U_g2513 (.A(G5014_2482_gat), .Y(G5018_2713_gat) );
OR5XL U_g2514 (.A(G4375_2521_gat), .B(G4374_2518_gat), .C(G4373_2519_gat), .D(G4372_2520_gat), .E(G4324_1284_gat), .Y(G4376_2714_gat) );
INVXL U_g2515 (.A(G4259_2487_gat), .Y(G4262_2715_gat) );
INVXL U_g2516 (.A(G4255_2488_gat), .Y(G4258_2716_gat) );
INVXL U_g2517 (.A(G3587_2489_gat), .Y(G3590_2717_gat) );
AND3XL U_g2518 (.A(G3591_2490_gat), .B(G3554_2510_gat), .C(G3563_2517_gat), .Y(G3611_2718_gat) );
INVXL U_g2519 (.A(G3591_2490_gat), .Y(G3594_2719_gat) );
OR4XL U_g2520 (.A(G4363_2465_gat), .B(G4362_2468_gat), .C(G4361_2470_gat), .D(G4297_1293_gat), .Y(G4364_2720_gat) );
OR2XL U_g2521 (.A(G89_48_ngat), .B(G4369_2486_ngat), .Y(G4380_2721_gat) );
INVXL U_g2522 (.A(G4614_2495_gat), .Y(G4617_2722_gat) );
AND3XL U_g2523 (.A(G4618_2496_gat), .B(G4581_2500_gat), .C(G4590_2499_gat), .Y(G4638_2723_gat) );
INVXL U_g2524 (.A(G4618_2496_gat), .Y(G4621_2724_gat) );
INVXL U_g2525 (.A(G3123_2497_gat), .Y(G3127_2725_gat) );
OR2XL U_g2526 (.A(G7617_2506_ngat), .B(G7614_2181_ngat), .Y(G7446_2726_gat) );
AND3XL U_g2527 (.A(G4614_2495_gat), .B(G4577_2183_gat), .C(G4586_2182_gat), .Y(G4635_2727_gat) );
INVXL U_g2528 (.A(G4610_2502_gat), .Y(G4613_2728_gat) );
INVXL U_g2529 (.A(G4606_2503_gat), .Y(G4609_2729_gat) );
AND3XL U_g2530 (.A(G4606_2503_gat), .B(G4554_1900_gat), .C(G4563_2184_gat), .Y(G4629_2730_gat) );
AND3XL U_g2531 (.A(G4610_2502_gat), .B(G4558_2189_gat), .C(G4567_2501_gat), .Y(G4632_2731_gat) );
OR2XL U_g2532 (.A(G6816_2515_ngat), .B(G6809_2190_ngat), .Y(G6818_2732_gat) );
OR4XL U_g2533 (.A(G3130_2513_gat), .B(G3129_2516_gat), .C(G3128_2509_gat), .D(G3059_1330_gat), .Y(G3131_2733_gat) );
OR2XL U_g2534 (.A(G6351_2505_ngat), .B(G6350_2514_ngat), .Y(G6352_2734_gat) );
OR2XL U_g2535 (.A(G7618_2498_ngat), .B(G7611_2193_ngat), .Y(G7447_2735_gat) );
OR2XL U_g2536 (.A(G7610_2508_ngat), .B(G7603_2196_ngat), .Y(G7457_2736_gat) );
OR2XL U_g2537 (.A(G7609_2507_ngat), .B(G7606_2197_ngat), .Y(G7456_2737_gat) );
OR5XL U_g2538 (.A(G3142_2478_gat), .B(G3141_2492_gat), .C(G3140_2494_gat), .D(G3139_2474_gat), .E(G3090_1356_gat), .Y(G3143_2738_gat) );
AND3XL U_g2539 (.A(G4255_2488_gat), .B(G4203_1923_gat), .C(G4212_1937_gat), .Y(G4278_2739_gat) );
AND3XL U_g2540 (.A(G4259_2487_gat), .B(G4207_2198_gat), .C(G4216_2206_gat), .Y(G4281_2740_gat) );
AND3XL U_g2541 (.A(G3587_2489_gat), .B(G3550_2199_gat), .C(G3559_2205_gat), .Y(G3608_2741_gat) );
INVXL U_g2542 (.A(G4980_2511_gat), .Y(G4986_2742_gat) );
INVXL U_g2543 (.A(G4939_2512_gat), .Y(G4945_2743_gat) );
OR2XL U_g2544 (.A(G6815_2504_ngat), .B(G6812_2204_ngat), .Y(G6817_2744_gat) );
BUFX20 U_g2545 (.A(G2472_2532_gat), .Y(G4836_2745_gat) );
BUFX20 U_g2546 (.A(G2742_2533_gat), .Y(G6294_2746_gat) );
BUFX20 U_g2547 (.A(G2742_2533_gat), .Y(G6206_2747_gat) );
AND3XL U_g2548 (.A(G1299_2536_gat), .B(G1253_2214_gat), .C(G1240_1950_gat), .Y(G1317_2748_gat) );
AND3XL U_g2549 (.A(G1295_2537_gat), .B(G1249_1952_gat), .C(G1244_2211_gat), .Y(G1314_2749_gat) );
OR2XL U_g2550 (.A(G6341_2538_ngat), .B(G6340_2539_ngat), .Y(G6342_2750_gat) );
OR2XL U_g2551 (.A(G5368_2541_ngat), .B(G5367_2540_ngat), .Y(G5388_2751_gat) );
AND3XL U_g2552 (.A(G1287_2544_gat), .B(G1226_1959_gat), .C(G1221_2222_gat), .Y(G1308_2752_gat) );
AND3XL U_g2553 (.A(G1291_2543_gat), .B(G1230_2221_gat), .C(G1217_1960_gat), .Y(G1311_2753_gat) );
OR2XL U_g2554 (.A(G4839_316_ngat), .B(G4836_2745_ngat), .Y(G371_2754_gat) );
OR2XL U_g2555 (.A(G4526_205_ngat), .B(G2771_2634_ngat), .Y(G2806_2755_gat) );
AND2XL U_g2556 (.A(G4526_205_gat), .B(G2508_2630_gat), .Y(G2563_2756_gat) );
AND2XL U_g2557 (.A(G4028_2579_gat), .B(G4004_2224_gat), .Y(G4090_2757_gat) );
OR2XL U_g2558 (.A(G6646_2556_ngat), .B(G6639_2560_ngat), .Y(G3470_2758_gat) );
OR2XL U_g2559 (.A(G6654_2557_ngat), .B(G6647_2559_ngat), .Y(G3473_2759_gat) );
AND2XL U_g2560 (.A(G3431_2229_gat), .B(G3453_2578_gat), .Y(G3467_2760_gat) );
INVXL U_g2561 (.A(G6647_2559_gat), .Y(G6653_2761_gat) );
INVXL U_g2562 (.A(G6639_2560_gat), .Y(G6645_2762_gat) );
INVXL U_g2563 (.A(G6996_2561_gat), .Y(G7000_2763_gat) );
INVXL U_g2564 (.A(G6938_2562_gat), .Y(G6942_2764_gat) );
OR2XL U_g2565 (.A(G6670_2563_ngat), .B(G6663_2567_ngat), .Y(G3480_2765_gat) );
OR2XL U_g2566 (.A(G6662_2564_ngat), .B(G6655_2568_ngat), .Y(G3477_2766_gat) );
INVXL U_g2567 (.A(G6663_2567_gat), .Y(G6669_2767_gat) );
INVXL U_g2568 (.A(G6655_2568_gat), .Y(G6661_2768_gat) );
INVXL U_g2569 (.A(G4017_2569_gat), .Y(G6986_2769_gat) );
OR2XL U_g2570 (.A(G4051_2247_gat), .B(G4017_2569_gat), .Y(G6928_2770_gat) );
OR2XL U_g2571 (.A(G6686_2570_ngat), .B(G6679_1469_ngat), .Y(G3488_2771_gat) );
OR2XL U_g2572 (.A(G6678_2571_ngat), .B(G6671_1116_ngat), .Y(G3484_2772_gat) );
INVXL U_g2573 (.A(G4028_2579_gat), .Y(G4032_2773_gat) );
INVXL U_g2574 (.A(G7152_2584_gat), .Y(G7156_2774_gat) );
INVXL U_g2575 (.A(G7064_2585_gat), .Y(G7068_2775_gat) );
INVXL U_g2576 (.A(G7132_2589_gat), .Y(G7136_2776_gat) );
INVXL U_g2577 (.A(G7044_2590_gat), .Y(G7048_2777_gat) );
INVXL U_g2578 (.A(G4048_2594_gat), .Y(G7142_2778_gat) );
OR2XL U_g2579 (.A(G4052_2292_gat), .B(G4048_2594_gat), .Y(G7054_2779_gat) );
OR2XL U_g2580 (.A(G7135_1780_ngat), .B(G7132_2589_ngat), .Y(G7137_2780_gat) );
OR2XL U_g2581 (.A(G7047_1485_ngat), .B(G7044_2590_ngat), .Y(G7049_2781_gat) );
INVXL U_g2582 (.A(G2495_2601_gat), .Y(G2499_2782_gat) );
INVXL U_g2583 (.A(G2757_2602_gat), .Y(G2761_2783_gat) );
AND2XL U_g2584 (.A(G2780_2629_gat), .B(G2749_2307_gat), .Y(G2853_2784_gat) );
AND2XL U_g2585 (.A(G2771_2634_gat), .B(G2749_2307_gat), .Y(G2852_2785_gat) );
OR2XL U_g2586 (.A(G5944_2606_ngat), .B(G5937_2610_ngat), .Y(G2542_2786_gat) );
OR2XL U_g2587 (.A(G5952_2607_ngat), .B(G5945_2609_ngat), .Y(G2545_2787_gat) );
AND2XL U_g2588 (.A(G2508_2630_gat), .B(G2487_2312_gat), .Y(G2532_2788_gat) );
AND2XL U_g2589 (.A(G2487_2312_gat), .B(G2515_2628_gat), .Y(G2536_2789_gat) );
INVXL U_g2590 (.A(G5945_2609_gat), .Y(G5951_2790_gat) );
INVXL U_g2591 (.A(G5937_2610_gat), .Y(G5943_2791_gat) );
INVXL U_g2592 (.A(G6128_2611_gat), .Y(G6132_2792_gat) );
INVXL U_g2593 (.A(G6070_2612_gat), .Y(G6074_2793_gat) );
OR2XL U_g2594 (.A(G5968_2613_ngat), .B(G5961_2617_ngat), .Y(G2552_2794_gat) );
OR2XL U_g2595 (.A(G5960_2614_ngat), .B(G5953_2618_ngat), .Y(G2549_2795_gat) );
INVXL U_g2596 (.A(G5961_2617_gat), .Y(G5967_2796_gat) );
INVXL U_g2597 (.A(G5953_2618_gat), .Y(G5959_2797_gat) );
INVXL U_g2598 (.A(G2768_2619_gat), .Y(G6118_2798_gat) );
OR2XL U_g2599 (.A(G2804_2327_gat), .B(G2768_2619_gat), .Y(G6060_2799_gat) );
OR2XL U_g2600 (.A(G5984_2622_ngat), .B(G5977_1493_ngat), .Y(G2560_2800_gat) );
OR2XL U_g2601 (.A(G5976_2623_ngat), .B(G5969_1137_ngat), .Y(G2556_2801_gat) );
INVXL U_g2602 (.A(G2780_2629_gat), .Y(G2784_2802_gat) );
INVXL U_g2603 (.A(G2771_2634_gat), .Y(G2775_2803_gat) );
OR5XL U_g2604 (.A(G2522_2550_gat), .B(G2520_2522_gat), .C(G2519_2361_gat), .D(G2518_2353_gat), .E(G2431_1140_gat), .Y(G4841_2804_gat) );
INVXL U_g2605 (.A(G6284_2635_gat), .Y(G6288_2805_gat) );
OR5XL U_g2606 (.A(G2791_2637_gat), .B(G2790_2526_gat), .C(G2789_2365_gat), .D(G2788_2356_gat), .E(G2670_1141_gat), .Y(G6196_2806_gat) );
OR4XL U_g2607 (.A(G2526_2549_gat), .B(G2524_2525_gat), .C(G2523_2363_gat), .D(G2448_1142_gat), .Y(G4849_2807_gat) );
INVXL U_g2608 (.A(G6264_2640_gat), .Y(G6268_2808_gat) );
OR4XL U_g2609 (.A(G2797_2644_gat), .B(G2796_2529_gat), .C(G2795_2368_gat), .D(G2693_1143_gat), .Y(G6176_2809_gat) );
OR3XL U_g2610 (.A(G2529_2548_gat), .B(G2527_2524_gat), .C(G2465_1144_gat), .Y(G4857_2810_gat) );
OR2XL U_g2611 (.A(G2807_2648_gat), .B(G2801_2645_gat), .Y(G6186_2811_gat) );
INVXL U_g2612 (.A(G2801_2645_gat), .Y(G6274_2812_gat) );
OR2XL U_g2613 (.A(G3045_2651_gat), .B(G3028_2372_gat), .Y(G3046_2813_gat) );
INVXL U_g2614 (.A(G7438_2650_gat), .Y(G7442_2814_gat) );
OR2XL U_g2615 (.A(G1789_2652_gat), .B(G1708_2378_gat), .Y(G1790_2815_gat) );
OR2XL U_g2616 (.A(G1981_2655_gat), .B(G1941_2379_gat), .Y(G1982_2816_gat) );
OR2XL U_g2617 (.A(G5823_2657_ngat), .B(G5820_2002_ngat), .Y(G1985_2817_gat) );
OR2XL U_g2618 (.A(G5831_2656_ngat), .B(G5828_2003_ngat), .Y(G1988_2818_gat) );
OR2XL U_g2619 (.A(G5847_2663_ngat), .B(G5844_2007_ngat), .Y(G1995_2819_gat) );
OR2XL U_g2620 (.A(G5839_2664_ngat), .B(G5836_2008_ngat), .Y(G1992_2820_gat) );
INVXL U_g2621 (.A(G5526_2662_gat), .Y(G5530_2821_gat) );
INVXL U_g2622 (.A(G5468_2665_gat), .Y(G5472_2822_gat) );
OR2XL U_g2623 (.A(G5529_1519_ngat), .B(G5526_2662_ngat), .Y(G5531_2823_gat) );
OR2XL U_g2624 (.A(G2004_2666_ngat), .B(G2003_2399_ngat), .Y(G2005_2824_gat) );
OR2XL U_g2625 (.A(G2000_2667_ngat), .B(G1999_2400_ngat), .Y(G2001_2825_gat) );
OR2XL U_g2626 (.A(G5471_1162_ngat), .B(G5468_2665_ngat), .Y(G5473_2826_gat) );
AND2XL U_g2627 (.A(G4626_2404_ngat), .B(G4625_2678_ngat), .Y(G4627_2827_gat) );
AND2XL U_g2628 (.A(G1721_2410_gat), .B(G1730_2668_gat), .Y(G1751_2828_gat) );
AND2XL U_g2629 (.A(G4623_2420_ngat), .B(G4622_2673_ngat), .Y(G4624_2829_gat) );
INVXL U_g2630 (.A(G5682_2674_gat), .Y(G5686_2830_gat) );
INVXL U_g2631 (.A(G5594_2675_gat), .Y(G5598_2831_gat) );
OR2XL U_g2632 (.A(G5676_2671_ngat), .B(G5669_1182_ngat), .Y(G5678_2832_gat) );
OR2XL U_g2633 (.A(G5588_2672_ngat), .B(G5581_911_ngat), .Y(G5590_2833_gat) );
OR2XL U_g2634 (.A(G4986_2742_ngat), .B(G4983_1191_ngat), .Y(G4988_2834_gat) );
OR2XL U_g2635 (.A(G1002_2682_gat), .B(G908_1192_gat), .Y(G265_2835_gat) );
OR2XL U_g2636 (.A(G4945_2743_ngat), .B(G4942_1551_ngat), .Y(G4947_2836_gat) );
OR2XL U_g2637 (.A(G1151_2681_gat), .B(G1117_1193_gat), .Y(G241_2837_gat) );
AND2XL U_g2638 (.A(G3599_2436_ngat), .B(G3598_2692_ngat), .Y(G3600_2838_gat) );
AND2XL U_g2639 (.A(G924_2441_gat), .B(G933_2683_gat), .Y(G962_2839_gat) );
INVXL U_g2640 (.A(G5112_2687_gat), .Y(G5116_2840_gat) );
AND2XL U_g2641 (.A(G3596_2450_ngat), .B(G3595_2688_ngat), .Y(G3597_2841_gat) );
INVXL U_g2642 (.A(G5024_2689_gat), .Y(G5028_2842_gat) );
OR2XL U_g2643 (.A(G5106_2712_ngat), .B(G5099_1218_ngat), .Y(G5108_2843_gat) );
OR2XL U_g2644 (.A(G5018_2713_ngat), .B(G5011_941_ngat), .Y(G5020_2844_gat) );
AND2XL U_g2645 (.A(G4284_2456_ngat), .B(G4283_2694_ngat), .Y(G4285_2845_gat) );
AND2XL U_g2646 (.A(G4287_2457_ngat), .B(G4286_2693_ngat), .Y(G4288_2846_gat) );
AND2XL U_g2647 (.A(G1321_2460_ngat), .B(G1320_2696_ngat), .Y(G1322_2847_gat) );
AND2XL U_g2648 (.A(G1324_2461_ngat), .B(G1323_2695_ngat), .Y(G1325_2848_gat) );
OR2XL U_g2649 (.A(G6361_2702_ngat), .B(G6360_2697_ngat), .Y(G6362_2849_gat) );
AND2XL U_g2650 (.A(G4376_2714_gat), .B(G4356_2466_gat), .Y(G4387_2850_gat) );
OR2XL U_g2651 (.A(G6828_2701_ngat), .B(G6827_2700_ngat), .Y(G6848_2851_gat) );
AND3XL U_g2652 (.A(G4254_2708_gat), .B(G4193_2493_gat), .C(G4180_2159_gat), .Y(G4274_2852_gat) );
AND3XL U_g2653 (.A(G3586_2704_gat), .B(G3540_2491_gat), .C(G3527_2160_gat), .Y(G3604_2853_gat) );
INVXL U_g2654 (.A(G4376_2714_gat), .Y(G4379_2854_gat) );
INVXL U_g2655 (.A(G4364_2720_gat), .Y(G4368_2855_gat) );
AND3XL U_g2656 (.A(G3582_2705_gat), .B(G3536_2174_gat), .C(G3531_2480_gat), .Y(G3601_2856_gat) );
AND3XL U_g2657 (.A(G4250_2709_gat), .B(G4189_2176_gat), .C(G4184_2479_gat), .Y(G4271_2857_gat) );
AND5XL U_g2658 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3156_2706_gat), .D(G4386_2698_gat), .E(G89_48_gat), .Y(G263_2858_gat) );
AND4XL U_g2659 (.A(G3035_2374_gat), .B(G3156_2706_gat), .C(G4386_2698_gat), .D(G89_48_gat), .Y(G3241_2859_gat) );
AND5XL U_g2660 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3156_2706_gat), .D(G4386_2698_gat), .E(G89_48_gat), .Y(G257_2860_gat) );
AND2XL U_g2661 (.A(G3143_2738_gat), .B(G3123_2497_gat), .Y(G3163_2861_gat) );
OR2XL U_g2662 (.A(G7447_2735_ngat), .B(G7446_2726_ngat), .Y(G7448_2862_gat) );
AND3XL U_g2663 (.A(G4617_2722_gat), .B(G4586_2182_gat), .C(G4581_2500_gat), .Y(G4634_2863_gat) );
AND3XL U_g2664 (.A(G4621_2724_gat), .B(G4590_2499_gat), .C(G4577_2183_gat), .Y(G4637_2864_gat) );
AND3XL U_g2665 (.A(G4609_2729_gat), .B(G4563_2184_gat), .C(G4558_2189_gat), .Y(G4628_2865_gat) );
AND3XL U_g2666 (.A(G4613_2728_gat), .B(G4567_2501_gat), .C(G4554_1900_gat), .Y(G4631_2866_gat) );
OR2XL U_g2667 (.A(G6818_2732_ngat), .B(G6817_2744_ngat), .Y(G6840_2867_gat) );
INVXL U_g2668 (.A(G3131_2733_gat), .Y(G3135_2868_gat) );
INVXL U_g2669 (.A(G6352_2734_gat), .Y(G6356_2869_gat) );
OR2XL U_g2670 (.A(G7457_2736_ngat), .B(G7456_2737_ngat), .Y(G7458_2870_gat) );
INVXL U_g2671 (.A(G3143_2738_gat), .Y(G3146_2871_gat) );
AND3XL U_g2672 (.A(G4262_2715_gat), .B(G4216_2206_gat), .C(G4203_1923_gat), .Y(G4280_2872_gat) );
AND3XL U_g2673 (.A(G3594_2719_gat), .B(G3563_2517_gat), .C(G3550_2199_gat), .Y(G3610_2873_gat) );
OR2XL U_g2674 (.A(G3258_2546_gat), .B(G3223_1698_gat), .Y(G3259_2874_gat) );
AND3XL U_g2675 (.A(G3590_2717_gat), .B(G3559_2205_gat), .C(G3554_2510_gat), .Y(G3607_2875_gat) );
AND3XL U_g2676 (.A(G4258_2716_gat), .B(G4212_1937_gat), .C(G4207_2198_gat), .Y(G4277_2876_gat) );
OR2XL U_g2677 (.A(G2531_2547_gat), .B(G2481_1721_gat), .Y(G4865_2877_gat) );
OR2XL U_g2678 (.A(G6267_2208_ngat), .B(G6264_2640_ngat), .Y(G6269_2878_gat) );
INVXL U_g2679 (.A(G4836_2745_gat), .Y(G4840_2879_gat) );
INVXL U_g2680 (.A(G6294_2746_gat), .Y(G6298_2880_gat) );
INVXL U_g2681 (.A(G6206_2747_gat), .Y(G6210_2881_gat) );
AND2XL U_g2682 (.A(G1315_2534_ngat), .B(G1314_2749_ngat), .Y(G1316_2882_gat) );
AND2XL U_g2683 (.A(G1318_2535_ngat), .B(G1317_2748_ngat), .Y(G1319_2883_gat) );
INVXL U_g2684 (.A(G6342_2750_gat), .Y(G6346_2884_gat) );
INVXL U_g2685 (.A(G5388_2751_gat), .Y(G5392_2885_gat) );
AND2XL U_g2686 (.A(G1312_2542_ngat), .B(G1311_2753_ngat), .Y(G1313_2886_gat) );
AND2XL U_g2687 (.A(G1309_2545_ngat), .B(G1308_2752_ngat), .Y(G1310_2887_gat) );
AND2XL U_g2688 (.A(G3249_2223_gat), .B(G3046_2813_gat), .Y(G254_2888_gat) );
AND2XL U_g2689 (.A(G3249_2223_gat), .B(G3046_2813_gat), .Y(G260_2889_gat) );
OR2XL U_g2690 (.A(G4840_2879_ngat), .B(G4833_207_ngat), .Y(G372_2890_gat) );
AND3XL U_g2691 (.A(G3466_2558_gat), .B(G2532_2788_gat), .C(G4526_205_gat), .Y(G3277_2891_gat) );
AND4XL U_g2692 (.A(G1974_2382_gat), .B(G3466_2558_gat), .C(G2532_2788_gat), .D(G4526_205_gat), .Y(G3270_2892_gat) );
AND2XL U_g2693 (.A(G2806_2755_gat), .B(G2784_2802_gat), .Y(G2809_2893_gat) );
AND3XL U_g2694 (.A(G4089_2553_gat), .B(G2852_2785_gat), .C(G4526_205_gat), .Y(G1454_2894_gat) );
AND4XL U_g2695 (.A(G1788_2375_gat), .B(G4089_2553_gat), .C(G2852_2785_gat), .D(G4526_205_gat), .Y(G1445_2895_gat) );
AND5XL U_g2696 (.A(G997_2432_gat), .B(G1788_2375_gat), .C(G4089_2553_gat), .D(G2852_2785_gat), .E(G4526_205_gat), .Y(G269_2896_gat) );
AND5XL U_g2697 (.A(G1146_2431_gat), .B(G1974_2382_gat), .C(G3466_2558_gat), .D(G2532_2788_gat), .E(G4526_205_gat), .Y(G245_2897_gat) );
OR2XL U_g2698 (.A(G3467_2760_gat), .B(G3437_2551_gat), .Y(G3468_2898_gat) );
OR2XL U_g2699 (.A(G4090_2757_gat), .B(G4010_2552_gat), .Y(G4091_2899_gat) );
OR2XL U_g2700 (.A(G6645_2762_ngat), .B(G6642_2227_ngat), .Y(G3469_2900_gat) );
OR2XL U_g2701 (.A(G6653_2761_ngat), .B(G6650_2228_ngat), .Y(G3472_2901_gat) );
OR2XL U_g2702 (.A(G6669_2767_ngat), .B(G6666_2232_ngat), .Y(G3479_2902_gat) );
OR2XL U_g2703 (.A(G6661_2768_ngat), .B(G6658_2233_ngat), .Y(G3476_2903_gat) );
INVXL U_g2704 (.A(G6986_2769_gat), .Y(G6990_2904_gat) );
INVXL U_g2705 (.A(G6928_2770_gat), .Y(G6932_2905_gat) );
OR2XL U_g2706 (.A(G3488_2771_ngat), .B(G3487_2574_ngat), .Y(G3489_2906_gat) );
OR2XL U_g2707 (.A(G6989_1769_ngat), .B(G6986_2769_ngat), .Y(G6991_2907_gat) );
OR2XL U_g2708 (.A(G6931_1471_ngat), .B(G6928_2770_ngat), .Y(G6933_2908_gat) );
OR2XL U_g2709 (.A(G3484_2772_ngat), .B(G3483_2577_ngat), .Y(G3485_2909_gat) );
AND2XL U_g2710 (.A(G4023_2582_gat), .B(G4032_2773_gat), .Y(G4053_2910_gat) );
INVXL U_g2711 (.A(G7142_2778_gat), .Y(G7146_2911_gat) );
INVXL U_g2712 (.A(G7054_2779_gat), .Y(G7058_2912_gat) );
OR2XL U_g2713 (.A(G7136_2776_ngat), .B(G7129_1483_ngat), .Y(G7138_2913_gat) );
OR2XL U_g2714 (.A(G7048_2777_ngat), .B(G7041_1127_ngat), .Y(G7050_2914_gat) );
OR2XL U_g2715 (.A(G2536_2789_gat), .B(G2495_2601_gat), .Y(G2537_2915_gat) );
OR2XL U_g2716 (.A(G2853_2784_gat), .B(G2757_2602_gat), .Y(G2854_2916_gat) );
OR2XL U_g2717 (.A(G2753_2603_ngat), .B(G2761_2783_ngat), .Y(G2808_2917_gat) );
OR2XL U_g2718 (.A(G5943_2791_ngat), .B(G5940_2310_ngat), .Y(G2541_2918_gat) );
OR2XL U_g2719 (.A(G5951_2790_ngat), .B(G5948_2311_ngat), .Y(G2544_2919_gat) );
OR2XL U_g2720 (.A(G2491_2608_ngat), .B(G2499_2782_ngat), .Y(G2577_2920_gat) );
OR2XL U_g2721 (.A(G5967_2796_ngat), .B(G5964_2315_ngat), .Y(G2551_2921_gat) );
OR2XL U_g2722 (.A(G5959_2797_ngat), .B(G5956_2316_ngat), .Y(G2548_2922_gat) );
INVXL U_g2723 (.A(G6118_2798_gat), .Y(G6122_2923_gat) );
INVXL U_g2724 (.A(G6060_2799_gat), .Y(G6064_2924_gat) );
OR2XL U_g2725 (.A(G2560_2800_ngat), .B(G2559_2624_ngat), .Y(G2561_2925_gat) );
OR2XL U_g2726 (.A(G6121_1790_ngat), .B(G6118_2798_ngat), .Y(G6123_2926_gat) );
OR2XL U_g2727 (.A(G6063_1495_ngat), .B(G6060_2799_ngat), .Y(G6065_2927_gat) );
OR2XL U_g2728 (.A(G2556_2801_ngat), .B(G2555_2627_ngat), .Y(G2557_2928_gat) );
OR2XL U_g2729 (.A(G2563_2756_gat), .B(G2515_2628_gat), .Y(G2564_2929_gat) );
AND2XL U_g2730 (.A(G2775_2803_gat), .B(G2784_2802_gat), .Y(G2813_2930_gat) );
OR2XL U_g2731 (.A(G4848_2631_ngat), .B(G4841_2804_ngat), .Y(G387_2931_gat) );
INVXL U_g2732 (.A(G4841_2804_gat), .Y(G4847_2932_gat) );
INVXL U_g2733 (.A(G6196_2806_gat), .Y(G6200_2933_gat) );
OR2XL U_g2734 (.A(G4856_2639_ngat), .B(G4849_2807_ngat), .Y(G390_2934_gat) );
INVXL U_g2735 (.A(G4849_2807_gat), .Y(G4855_2935_gat) );
INVXL U_g2736 (.A(G6176_2809_gat), .Y(G6180_2936_gat) );
OR2XL U_g2737 (.A(G4864_2641_ngat), .B(G4857_2810_ngat), .Y(G393_2937_gat) );
INVXL U_g2738 (.A(G4857_2810_gat), .Y(G4863_2938_gat) );
INVXL U_g2739 (.A(G6186_2811_gat), .Y(G6190_2939_gat) );
INVXL U_g2740 (.A(G6274_2812_gat), .Y(G6278_2940_gat) );
OR2XL U_g2741 (.A(G4872_2649_ngat), .B(G4865_2877_ngat), .Y(G396_2941_gat) );
OR2XL U_g2742 (.A(G1986_2653_ngat), .B(G1985_2817_ngat), .Y(G1987_2942_gat) );
OR2XL U_g2743 (.A(G1989_2654_ngat), .B(G1988_2818_ngat), .Y(G1990_2943_gat) );
OR2XL U_g2744 (.A(G1996_2658_ngat), .B(G1995_2819_ngat), .Y(G1997_2944_gat) );
OR2XL U_g2745 (.A(G1993_2659_ngat), .B(G1992_2820_ngat), .Y(G1994_2945_gat) );
OR2XL U_g2746 (.A(G5530_2821_ngat), .B(G5523_1158_ngat), .Y(G5532_2946_gat) );
INVXL U_g2747 (.A(G2001_2825_gat), .Y(G2002_2947_gat) );
OR2XL U_g2748 (.A(G5472_2822_ngat), .B(G5465_885_ngat), .Y(G5474_2948_gat) );
OR2XL U_g2749 (.A(G4624_2829_ngat), .B(G4627_2827_ngat), .Y(G7433_2949_gat) );
INVXL U_g2750 (.A(G1751_2828_gat), .Y(G1754_2950_gat) );
OR2XL U_g2751 (.A(G5678_2832_ngat), .B(G5677_2676_ngat), .Y(G5679_2951_gat) );
OR2XL U_g2752 (.A(G5590_2833_ngat), .B(G5589_2677_ngat), .Y(G5591_2952_gat) );
OR2XL U_g2753 (.A(G4989_2679_ngat), .B(G4988_2834_ngat), .Y(G4990_2953_gat) );
OR2XL U_g2754 (.A(G4948_2680_ngat), .B(G4947_2836_ngat), .Y(G4949_2954_gat) );
AND2XL U_g2755 (.A(G1146_2431_gat), .B(G1982_2816_gat), .Y(G242_2955_gat) );
AND2XL U_g2756 (.A(G997_2432_gat), .B(G1790_2815_gat), .Y(G266_2956_gat) );
OR2XL U_g2757 (.A(G3597_2841_ngat), .B(G3600_2838_ngat), .Y(G6829_2957_gat) );
INVXL U_g2758 (.A(G962_2839_gat), .Y(G965_2958_gat) );
OR2XL U_g2759 (.A(G5108_2843_ngat), .B(G5107_2690_ngat), .Y(G5109_2959_gat) );
OR2XL U_g2760 (.A(G5020_2844_ngat), .B(G5019_2691_ngat), .Y(G5021_2960_gat) );
OR2XL U_g2761 (.A(G4285_2845_ngat), .B(G4288_2846_ngat), .Y(G6337_2961_gat) );
OR2XL U_g2762 (.A(G1322_2847_ngat), .B(G1325_2848_ngat), .Y(G5385_2962_gat) );
INVXL U_g2763 (.A(G6362_2849_gat), .Y(G6366_2963_gat) );
OR2XL U_g2764 (.A(G4360_2699_ngat), .B(G4368_2855_ngat), .Y(G4381_2964_gat) );
INVXL U_g2765 (.A(G6848_2851_gat), .Y(G6852_2965_gat) );
AND2XL U_g2766 (.A(G3605_2703_ngat), .B(G3604_2853_ngat), .Y(G3606_2966_gat) );
AND2XL U_g2767 (.A(G4275_2707_ngat), .B(G4274_2852_ngat), .Y(G4276_2967_gat) );
AND2XL U_g2768 (.A(G4272_2710_ngat), .B(G4271_2857_ngat), .Y(G4273_2968_gat) );
AND2XL U_g2769 (.A(G3602_2711_ngat), .B(G3601_2856_ngat), .Y(G3603_2969_gat) );
AND2XL U_g2770 (.A(G3611_2718_ngat), .B(G3610_2873_ngat), .Y(G3612_2970_gat) );
OR2XL U_g2771 (.A(G4387_2850_gat), .B(G4364_2720_gat), .Y(G4388_2971_gat) );
AND2XL U_g2772 (.A(G4380_2721_gat), .B(G4379_2854_gat), .Y(G4382_2972_gat) );
AND2XL U_g2773 (.A(G4638_2723_ngat), .B(G4637_2864_ngat), .Y(G4639_2973_gat) );
OR2XL U_g2774 (.A(G3127_2725_ngat), .B(G3135_2868_ngat), .Y(G3151_2974_gat) );
INVXL U_g2775 (.A(G7448_2862_gat), .Y(G7452_2975_gat) );
AND2XL U_g2776 (.A(G4635_2727_ngat), .B(G4634_2863_ngat), .Y(G4636_2976_gat) );
AND2XL U_g2777 (.A(G4629_2730_ngat), .B(G4628_2865_ngat), .Y(G4630_2977_gat) );
AND2XL U_g2778 (.A(G4632_2731_ngat), .B(G4631_2866_ngat), .Y(G4633_2978_gat) );
INVXL U_g2779 (.A(G6840_2867_gat), .Y(G6844_2979_gat) );
OR2XL U_g2780 (.A(G3163_2861_gat), .B(G3131_2733_gat), .Y(G3164_2980_gat) );
INVXL U_g2781 (.A(G7458_2870_gat), .Y(G7462_2981_gat) );
AND2XL U_g2782 (.A(G4278_2739_ngat), .B(G4277_2876_ngat), .Y(G4279_2982_gat) );
AND2XL U_g2783 (.A(G4281_2740_ngat), .B(G4280_2872_ngat), .Y(G4282_2983_gat) );
AND2XL U_g2784 (.A(G3608_2741_ngat), .B(G3607_2875_ngat), .Y(G3609_2984_gat) );
INVXL U_g2785 (.A(G4865_2877_gat), .Y(G4871_2985_gat) );
OR2XL U_g2786 (.A(G6268_2808_ngat), .B(G6261_1944_ngat), .Y(G6270_2986_gat) );
OR2XL U_g2787 (.A(G6179_1946_ngat), .B(G6176_2809_ngat), .Y(G6181_2987_gat) );
OR2XL U_g2788 (.A(G1316_2882_ngat), .B(G1319_2883_ngat), .Y(G5377_2988_gat) );
OR2XL U_g2789 (.A(G1310_2887_ngat), .B(G1313_2886_ngat), .Y(G5369_2989_gat) );
AND3XL U_g2790 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3164_2980_gat), .Y(G255_2990_gat) );
AND4XL U_g2791 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3156_2706_gat), .D(G4388_2971_gat), .Y(G256_2991_gat) );
AND3XL U_g2792 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3164_2980_gat), .Y(G261_2992_gat) );
AND4XL U_g2793 (.A(G3249_2223_gat), .B(G3035_2374_gat), .C(G3156_2706_gat), .D(G4388_2971_gat), .Y(G262_2993_gat) );
INVXL U_g2794 (.A(G2809_2893_gat), .Y(G2812_2995_gat) );
AND2XL U_g2795 (.A(G4089_2553_gat), .B(G2854_2916_gat), .Y(G1450_2996_gat) );
OR2XL U_g2796 (.A(G3470_2758_ngat), .B(G3469_2900_ngat), .Y(G3471_2997_gat) );
OR2XL U_g2797 (.A(G3473_2759_ngat), .B(G3472_2901_ngat), .Y(G3474_2998_gat) );
AND2XL U_g2798 (.A(G3466_2558_gat), .B(G2537_2915_gat), .Y(G3274_2999_gat) );
OR2XL U_g2799 (.A(G3480_2765_ngat), .B(G3479_2902_ngat), .Y(G3481_3000_gat) );
OR2XL U_g2800 (.A(G3477_2766_ngat), .B(G3476_2903_ngat), .Y(G3478_3001_gat) );
OR2XL U_g2801 (.A(G6990_2904_ngat), .B(G6983_1470_ngat), .Y(G6992_3002_gat) );
OR2XL U_g2802 (.A(G6932_2905_ngat), .B(G6925_1115_ngat), .Y(G6934_3003_gat) );
INVXL U_g2803 (.A(G3485_2909_gat), .Y(G3486_3004_gat) );
INVXL U_g2804 (.A(G4053_2910_gat), .Y(G4056_3005_gat) );
OR2XL U_g2805 (.A(G7138_2913_ngat), .B(G7137_2780_ngat), .Y(G7139_3006_gat) );
OR2XL U_g2806 (.A(G7050_2914_ngat), .B(G7049_2781_ngat), .Y(G7051_3007_gat) );
AND2XL U_g2807 (.A(G2757_2602_gat), .B(G2809_2893_gat), .Y(G2851_3008_gat) );
OR2XL U_g2808 (.A(G2542_2786_ngat), .B(G2541_2918_ngat), .Y(G2543_3009_gat) );
OR2XL U_g2809 (.A(G2545_2787_ngat), .B(G2544_2919_ngat), .Y(G2546_3010_gat) );
AND2XL U_g2810 (.A(G2564_2929_gat), .B(G2577_2920_gat), .Y(G2579_3011_gat) );
OR2XL U_g2811 (.A(G2552_2794_ngat), .B(G2551_2921_ngat), .Y(G2553_3012_gat) );
OR2XL U_g2812 (.A(G2549_2795_ngat), .B(G2548_2922_ngat), .Y(G2550_3013_gat) );
OR2XL U_g2813 (.A(G6122_2923_ngat), .B(G6115_1494_ngat), .Y(G6124_3014_gat) );
OR2XL U_g2814 (.A(G6064_2924_ngat), .B(G6057_1136_ngat), .Y(G6066_3015_gat) );
AND2XL U_g2815 (.A(G2406_2344_gat), .B(G2564_2929_gat), .Y(G384_3016_gat) );
INVXL U_g2816 (.A(G2557_2928_gat), .Y(G2558_3017_gat) );
INVXL U_g2817 (.A(G2564_2929_gat), .Y(G2571_3018_gat) );
INVXL U_g2818 (.A(G2813_2930_gat), .Y(G2816_3019_gat) );
OR2XL U_g2819 (.A(G4847_2932_ngat), .B(G4844_2345_ngat), .Y(G386_3020_gat) );
OR2XL U_g2820 (.A(G4855_2935_ngat), .B(G4852_2352_ngat), .Y(G389_3021_gat) );
OR2XL U_g2821 (.A(G4863_2938_ngat), .B(G4860_2358_ngat), .Y(G392_3022_gat) );
OR2XL U_g2822 (.A(G4871_2985_ngat), .B(G4868_2371_ngat), .Y(G395_3023_gat) );
OR2XL U_g2823 (.A(G7442_2814_ngat), .B(G7433_2949_ngat), .Y(G4516_3024_gat) );
AND2XL U_g2824 (.A(G3035_2374_gat), .B(G3164_2980_gat), .Y(G3239_3025_gat) );
AND3XL U_g2825 (.A(G3035_2374_gat), .B(G3156_2706_gat), .C(G4388_2971_gat), .Y(G3240_3026_gat) );
AND3XL U_g2826 (.A(G997_2432_gat), .B(G1788_2375_gat), .C(G4091_2899_gat), .Y(G267_3027_gat) );
AND4XL U_g2827 (.A(G997_2432_gat), .B(G1788_2375_gat), .C(G4089_2553_gat), .D(G2854_2916_gat), .Y(G268_3028_gat) );
AND2XL U_g2828 (.A(G1788_2375_gat), .B(G4091_2899_gat), .Y(G1436_3029_gat) );
AND3XL U_g2829 (.A(G1788_2375_gat), .B(G4089_2553_gat), .C(G2854_2916_gat), .Y(G1440_3030_gat) );
INVXL U_g2830 (.A(G1990_2943_gat), .Y(G1991_3031_gat) );
AND3XL U_g2831 (.A(G1146_2431_gat), .B(G1974_2382_gat), .C(G3468_2898_gat), .Y(G243_3032_gat) );
AND4XL U_g2832 (.A(G1146_2431_gat), .B(G1974_2382_gat), .C(G3466_2558_gat), .D(G2537_2915_gat), .Y(G244_3033_gat) );
AND2XL U_g2833 (.A(G1974_2382_gat), .B(G3468_2898_gat), .Y(G3265_3034_gat) );
AND3XL U_g2834 (.A(G1974_2382_gat), .B(G3466_2558_gat), .C(G2537_2915_gat), .Y(G3267_3035_gat) );
INVXL U_g2835 (.A(G1997_2944_gat), .Y(G1998_3036_gat) );
OR2XL U_g2836 (.A(G5532_2946_ngat), .B(G5531_2823_ngat), .Y(G5533_3037_gat) );
OR2XL U_g2837 (.A(G5474_2948_ngat), .B(G5473_2826_ngat), .Y(G5475_3038_gat) );
INVXL U_g2838 (.A(G7433_2949_gat), .Y(G7441_3039_gat) );
OR2XL U_g2839 (.A(G5686_2830_ngat), .B(G5679_2951_ngat), .Y(G5688_3040_gat) );
OR2XL U_g2840 (.A(G5598_2831_ngat), .B(G5591_2952_ngat), .Y(G5600_3041_gat) );
INVXL U_g2841 (.A(G5679_2951_gat), .Y(G5685_3042_gat) );
INVXL U_g2842 (.A(G5591_2952_gat), .Y(G5597_3043_gat) );
OR2XL U_g2843 (.A(G6836_1833_ngat), .B(G6829_2957_ngat), .Y(G3614_3044_gat) );
INVXL U_g2844 (.A(G4990_2953_gat), .Y(G4996_3045_gat) );
INVXL U_g2845 (.A(G4949_2954_gat), .Y(G4955_3046_gat) );
OR2XL U_g2846 (.A(G4997_1555_ngat), .B(G4990_2953_ngat), .Y(G4999_3047_gat) );
OR2XL U_g2847 (.A(G4956_1556_ngat), .B(G4949_2954_ngat), .Y(G4958_3048_gat) );
INVXL U_g2848 (.A(G6829_2957_gat), .Y(G6835_3049_gat) );
OR2XL U_g2849 (.A(G5116_2840_ngat), .B(G5109_2959_ngat), .Y(G5118_3050_gat) );
OR2XL U_g2850 (.A(G5028_2842_ngat), .B(G5021_2960_ngat), .Y(G5030_3051_gat) );
INVXL U_g2851 (.A(G5109_2959_gat), .Y(G5115_3052_gat) );
INVXL U_g2852 (.A(G5021_2960_gat), .Y(G5027_3053_gat) );
INVXL U_g2853 (.A(G6337_2961_gat), .Y(G6345_3054_gat) );
INVXL U_g2854 (.A(G5385_2962_gat), .Y(G5391_3055_gat) );
OR2XL U_g2855 (.A(G3603_2969_ngat), .B(G3606_2966_ngat), .Y(G6837_3056_gat) );
OR2XL U_g2856 (.A(G4273_2968_ngat), .B(G4276_2967_ngat), .Y(G6347_3057_gat) );
OR2XL U_g2857 (.A(G3609_2984_ngat), .B(G3612_2970_ngat), .Y(G6845_3058_gat) );
AND2XL U_g2858 (.A(G4364_2720_gat), .B(G4382_2972_gat), .Y(G3148_3059_gat) );
INVXL U_g2859 (.A(G4382_2972_gat), .Y(G4385_3060_gat) );
OR2XL U_g2860 (.A(G4636_2976_ngat), .B(G4639_2973_ngat), .Y(G7443_3061_gat) );
OR2XL U_g2861 (.A(G4630_2977_ngat), .B(G4633_2978_ngat), .Y(G7453_3062_gat) );
OR2XL U_g2862 (.A(G4279_2982_ngat), .B(G4282_2983_ngat), .Y(G6357_3063_gat) );
OR2XL U_g2863 (.A(G6270_2986_ngat), .B(G6269_2878_ngat), .Y(G6271_3064_gat) );
OR2XL U_g2864 (.A(G6180_2936_ngat), .B(G6173_1723_ngat), .Y(G6182_3065_gat) );
INVXL U_g2865 (.A(G5377_2988_gat), .Y(G5383_3066_gat) );
OR2XL U_g2866 (.A(G5384_1953_ngat), .B(G5377_2988_ngat), .Y(G1330_3067_gat) );
OR2XL U_g2867 (.A(G6346_2884_ngat), .B(G6337_2961_ngat), .Y(G2860_3068_gat) );
OR2XL U_g2868 (.A(G5392_2885_ngat), .B(G5385_2962_ngat), .Y(G1333_3069_gat) );
INVXL U_g2869 (.A(G5369_2989_gat), .Y(G5375_3070_gat) );
OR2XL U_g2870 (.A(G5376_1961_ngat), .B(G5369_2989_ngat), .Y(G1327_3071_gat) );
OR3XL U_g2871 (.A(G3277_2891_gat), .B(G3274_2999_gat), .C(G3468_2898_gat), .Y(G3279_3072_gat) );
OR3XL U_g2872 (.A(G1454_2894_gat), .B(G1450_2996_gat), .C(G4091_2899_gat), .Y(G1766_3073_gat) );
INVXL U_g2873 (.A(G3474_2998_gat), .Y(G3475_3074_gat) );
INVXL U_g2874 (.A(G3481_3000_gat), .Y(G3482_3075_gat) );
OR2XL U_g2875 (.A(G6992_3002_ngat), .B(G6991_2907_ngat), .Y(G6993_3076_gat) );
OR2XL U_g2876 (.A(G6934_3003_ngat), .B(G6933_2908_ngat), .Y(G6935_3077_gat) );
OR2XL U_g2877 (.A(G7146_2911_ngat), .B(G7139_3006_ngat), .Y(G7148_3078_gat) );
OR2XL U_g2878 (.A(G7058_2912_ngat), .B(G7051_3007_ngat), .Y(G7060_3079_gat) );
INVXL U_g2879 (.A(G7139_3006_gat), .Y(G7145_3080_gat) );
INVXL U_g2880 (.A(G7051_3007_gat), .Y(G7057_3081_gat) );
AND2XL U_g2881 (.A(G2571_3018_gat), .B(G2495_2601_gat), .Y(G2578_3082_gat) );
AND2XL U_g2882 (.A(G2812_2995_gat), .B(G2808_2917_gat), .Y(G2850_3083_gat) );
INVXL U_g2883 (.A(G2546_3010_gat), .Y(G2547_3084_gat) );
INVXL U_g2884 (.A(G2553_3012_gat), .Y(G2554_3085_gat) );
AND2XL U_g2885 (.A(G2571_3018_gat), .B(G2561_2925_gat), .Y(G380_3086_gat) );
OR2XL U_g2886 (.A(G6124_3014_ngat), .B(G6123_2926_ngat), .Y(G6125_3087_gat) );
OR2XL U_g2887 (.A(G6066_3015_ngat), .B(G6065_2927_ngat), .Y(G6067_3088_gat) );
AND2XL U_g2888 (.A(G2571_3018_gat), .B(G2400_1988_gat), .Y(G383_3089_gat) );
AND2XL U_g2889 (.A(G2543_3009_gat), .B(G2564_2929_gat), .Y(G375_3090_gat) );
AND2XL U_g2890 (.A(G2550_3013_gat), .B(G2564_2929_gat), .Y(G378_3091_gat) );
AND2XL U_g2891 (.A(G2558_3017_gat), .B(G2564_2929_gat), .Y(G381_3092_gat) );
OR2XL U_g2892 (.A(G6278_2940_ngat), .B(G6271_3064_ngat), .Y(G6280_3096_gat) );
OR4XL U_g2893 (.A(G3241_2859_gat), .B(G3240_3026_gat), .C(G3239_3025_gat), .D(G3046_2813_gat), .Y(G3242_3098_gat) );
OR2XL U_g2894 (.A(G7441_3039_ngat), .B(G7438_2650_ngat), .Y(G4515_3099_gat) );
OR4XL U_g2895 (.A(G1445_2895_gat), .B(G1440_3030_gat), .C(G1436_3029_gat), .D(G1790_2815_gat), .Y(G1447_3100_gat) );
OR4XL U_g2896 (.A(G3270_2892_gat), .B(G3267_3035_gat), .C(G3265_3034_gat), .D(G1982_2816_gat), .Y(G3271_3101_gat) );
OR2XL U_g2897 (.A(G5540_2660_ngat), .B(G5533_3037_ngat), .Y(G5542_3102_gat) );
OR2XL U_g2898 (.A(G5482_2661_ngat), .B(G5475_3038_ngat), .Y(G5484_3103_gat) );
INVXL U_g2899 (.A(G5533_3037_gat), .Y(G5539_3104_gat) );
INVXL U_g2900 (.A(G5475_3038_gat), .Y(G5481_3105_gat) );
OR2XL U_g2901 (.A(G5685_3042_ngat), .B(G5682_2674_ngat), .Y(G5687_3106_gat) );
OR2XL U_g2902 (.A(G5597_3043_ngat), .B(G5594_2675_ngat), .Y(G5599_3107_gat) );
OR2XL U_g2903 (.A(G6835_3049_ngat), .B(G6832_1546_ngat), .Y(G3613_3108_gat) );
OR2XL U_g2904 (.A(G4996_3045_ngat), .B(G4993_1203_ngat), .Y(G4998_3111_gat) );
OR2XL U_g2905 (.A(G4955_3046_ngat), .B(G4952_1204_ngat), .Y(G4957_3112_gat) );
OR2XL U_g2906 (.A(G5115_3052_ngat), .B(G5112_2687_ngat), .Y(G5117_3113_gat) );
OR2XL U_g2907 (.A(G5027_3053_ngat), .B(G5024_2689_ngat), .Y(G5029_3114_gat) );
OR2XL U_g2908 (.A(G6366_2963_ngat), .B(G6357_3063_ngat), .Y(G2866_3115_gat) );
AND2XL U_g2909 (.A(G4385_3060_gat), .B(G4381_2964_gat), .Y(G3147_3116_gat) );
OR2XL U_g2910 (.A(G6852_2965_ngat), .B(G6845_3058_ngat), .Y(G3620_3117_gat) );
INVXL U_g2911 (.A(G6837_3056_gat), .Y(G6843_3118_gat) );
INVXL U_g2912 (.A(G6347_3057_gat), .Y(G6355_3119_gat) );
INVXL U_g2913 (.A(G6845_3058_gat), .Y(G6851_3120_gat) );
INVXL U_g2914 (.A(G7443_3061_gat), .Y(G7451_3123_gat) );
OR2XL U_g2915 (.A(G7452_2975_ngat), .B(G7443_3061_ngat), .Y(G4519_3124_gat) );
INVXL U_g2916 (.A(G7453_3062_gat), .Y(G7461_3125_gat) );
OR2XL U_g2917 (.A(G6844_2979_ngat), .B(G6837_3056_ngat), .Y(G3617_3126_gat) );
OR2XL U_g2918 (.A(G6356_2869_ngat), .B(G6347_3057_ngat), .Y(G2863_3127_gat) );
OR2XL U_g2919 (.A(G7462_2981_ngat), .B(G7453_3062_ngat), .Y(G4522_3128_gat) );
INVXL U_g2920 (.A(G6357_3063_gat), .Y(G6365_3129_gat) );
INVXL U_g2921 (.A(G6271_3064_gat), .Y(G6277_3130_gat) );
OR2XL U_g2922 (.A(G6182_3065_ngat), .B(G6181_2987_ngat), .Y(G6183_3131_gat) );
OR2XL U_g2923 (.A(G5383_3066_ngat), .B(G5380_1736_ngat), .Y(G1329_3132_gat) );
OR2XL U_g2924 (.A(G6345_3054_ngat), .B(G6342_2750_ngat), .Y(G2859_3133_gat) );
OR2XL U_g2925 (.A(G5391_3055_ngat), .B(G5388_2751_ngat), .Y(G1332_3134_gat) );
OR2XL U_g2926 (.A(G5375_3070_ngat), .B(G5372_1759_ngat), .Y(G1326_3135_gat) );
BUFX20 U_g2927 (.A(G3279_3072_gat), .Y(G4713_3136_gat) );
INVXL U_g2928 (.A(G1766_3073_gat), .Y(G1771_3137_gat) );
OR2XL U_g2929 (.A(G7000_2763_ngat), .B(G6993_3076_ngat), .Y(G7002_3138_gat) );
OR2XL U_g2930 (.A(G6942_2764_ngat), .B(G6935_3077_ngat), .Y(G6944_3139_gat) );
INVXL U_g2931 (.A(G6993_3076_gat), .Y(G6999_3140_gat) );
INVXL U_g2932 (.A(G6935_3077_gat), .Y(G6941_3141_gat) );
OR2XL U_g2933 (.A(G7145_3080_ngat), .B(G7142_2778_ngat), .Y(G7147_3142_gat) );
OR2XL U_g2934 (.A(G7057_3081_ngat), .B(G7054_2779_ngat), .Y(G7059_3143_gat) );
OR2XL U_g2935 (.A(G2851_3008_gat), .B(G2850_3083_gat), .Y(G4067_3144_gat) );
OR2XL U_g2936 (.A(G2579_3011_gat), .B(G2578_3082_gat), .Y(G2580_3145_gat) );
OR2XL U_g2937 (.A(G6132_2792_ngat), .B(G6125_3087_ngat), .Y(G6134_3146_gat) );
OR2XL U_g2938 (.A(G6074_2793_ngat), .B(G6067_3088_ngat), .Y(G6076_3147_gat) );
INVXL U_g2939 (.A(G6125_3087_gat), .Y(G6131_3149_gat) );
INVXL U_g2940 (.A(G6067_3088_gat), .Y(G6073_3150_gat) );
AND2XL U_g2941 (.A(G2571_3018_gat), .B(G2547_3084_gat), .Y(G374_3152_gat) );
AND2XL U_g2942 (.A(G2571_3018_gat), .B(G2554_3085_gat), .Y(G377_3153_gat) );
OR2XL U_g2943 (.A(G6190_2939_ngat), .B(G6183_3131_ngat), .Y(G6192_3154_gat) );
OR2XL U_g2944 (.A(G6277_3130_ngat), .B(G6274_2812_ngat), .Y(G6279_3155_gat) );
OR2XL U_g2945 (.A(G4516_3024_ngat), .B(G4515_3099_ngat), .Y(G4517_3156_gat) );
BUFX20 U_g2946 (.A(G1447_3100_gat), .Y(G975_3157_gat) );
BUFX20 U_g2947 (.A(G3271_3101_gat), .Y(G4753_3158_gat) );
OR2XL U_g2948 (.A(G5539_3104_ngat), .B(G5536_2387_ngat), .Y(G5541_3159_gat) );
OR2XL U_g2949 (.A(G5481_3105_ngat), .B(G5478_2388_ngat), .Y(G5483_3160_gat) );
AND2XL U_g2950 (.A(G3279_3072_gat), .B(G1950_2047_gat), .Y(G2007_3161_gat) );
AND5XL U_g2951 (.A(G1869_1819_gat), .B(G1903_1826_gat), .C(G1885_1825_gat), .D(G1921_1832_gat), .E(G3279_3072_gat), .Y(G1964_3162_gat) );
AND4XL U_g2952 (.A(G1903_1826_gat), .B(G1885_1825_gat), .C(G1921_1832_gat), .D(G3279_3072_gat), .Y(G1968_3163_gat) );
OR2XL U_g2953 (.A(G5688_3040_ngat), .B(G5687_3106_ngat), .Y(G5689_3164_gat) );
AND3XL U_g2954 (.A(G1903_1826_gat), .B(G1921_1832_gat), .C(G3279_3072_gat), .Y(G1971_3165_gat) );
OR2XL U_g2955 (.A(G5600_3041_ngat), .B(G5599_3107_ngat), .Y(G5601_3166_gat) );
AND2XL U_g2956 (.A(G1921_1832_gat), .B(G3279_3072_gat), .Y(G1973_3167_gat) );
OR2XL U_g2957 (.A(G3614_3044_ngat), .B(G3613_3108_ngat), .Y(G3615_3168_gat) );
OR2XL U_g2958 (.A(G4999_3047_ngat), .B(G4998_3111_ngat), .Y(G5000_3169_gat) );
OR2XL U_g2959 (.A(G4958_3048_ngat), .B(G4957_3112_ngat), .Y(G4959_3170_gat) );
OR2XL U_g2960 (.A(G3242_3098_ngat), .B(G3228_2097_ngat), .Y(G3243_3171_gat) );
OR2XL U_g2961 (.A(G1447_3100_ngat), .B(G920_2100_ngat), .Y(G955_3172_gat) );
AND2XL U_g2962 (.A(G3271_3101_gat), .B(G1122_2101_gat), .Y(G1160_3173_gat) );
AND5XL U_g2963 (.A(G1038_1843_gat), .B(G1074_1846_gat), .C(G1055_1875_gat), .D(G1093_1853_gat), .E(G3271_3101_gat), .Y(G1136_3174_gat) );
OR2XL U_g2964 (.A(G5118_3050_ngat), .B(G5117_3113_ngat), .Y(G5119_3175_gat) );
AND4XL U_g2965 (.A(G1074_1846_gat), .B(G1055_1875_gat), .C(G1093_1853_gat), .D(G3271_3101_gat), .Y(G1140_3176_gat) );
AND3XL U_g2966 (.A(G1074_1846_gat), .B(G1093_1853_gat), .C(G3271_3101_gat), .Y(G1143_3177_gat) );
OR2XL U_g2967 (.A(G5030_3051_ngat), .B(G5029_3114_ngat), .Y(G5031_3178_gat) );
AND2XL U_g2968 (.A(G1093_1853_gat), .B(G3271_3101_gat), .Y(G1145_3179_gat) );
OR2XL U_g2969 (.A(G6365_3129_ngat), .B(G6362_2849_ngat), .Y(G2865_3180_gat) );
OR2XL U_g2970 (.A(G6851_3120_ngat), .B(G6848_2851_ngat), .Y(G3619_3181_gat) );
OR2XL U_g2971 (.A(G3148_3059_gat), .B(G3147_3116_gat), .Y(G3149_3182_gat) );
OR2XL U_g2972 (.A(G7451_3123_ngat), .B(G7448_2862_ngat), .Y(G4518_3183_gat) );
OR2XL U_g2973 (.A(G6843_3118_ngat), .B(G6840_2867_ngat), .Y(G3616_3184_gat) );
OR2XL U_g2974 (.A(G6355_3119_ngat), .B(G6352_2734_ngat), .Y(G2862_3185_gat) );
OR2XL U_g2975 (.A(G7461_3125_ngat), .B(G7458_2870_ngat), .Y(G4521_3186_gat) );
INVXL U_g2976 (.A(G6183_3131_gat), .Y(G6189_3187_gat) );
OR2XL U_g2977 (.A(G1330_3067_ngat), .B(G1329_3132_ngat), .Y(G1331_3188_gat) );
OR2XL U_g2978 (.A(G2860_3068_ngat), .B(G2859_3133_ngat), .Y(G2861_3189_gat) );
OR2XL U_g2979 (.A(G1333_3069_ngat), .B(G1332_3134_ngat), .Y(G1334_3190_gat) );
OR2XL U_g2980 (.A(G1327_3071_ngat), .B(G1326_3135_ngat), .Y(G1328_3191_gat) );
INVXL U_g2981 (.A(G4713_3136_gat), .Y(G4719_3192_gat) );
OR2XL U_g2982 (.A(G6999_3140_ngat), .B(G6996_2561_ngat), .Y(G7001_3193_gat) );
OR2XL U_g2983 (.A(G6941_3141_ngat), .B(G6938_2562_ngat), .Y(G6943_3194_gat) );
AND2XL U_g2984 (.A(G2580_3145_gat), .B(G3446_2265_gat), .Y(G3490_3195_gat) );
AND5XL U_g2985 (.A(G3365_1973_gat), .B(G3399_1978_gat), .C(G3381_1976_gat), .D(G3417_1979_gat), .E(G2580_3145_gat), .Y(G3459_3196_gat) );
AND4XL U_g2986 (.A(G3399_1978_gat), .B(G3381_1976_gat), .C(G3417_1979_gat), .D(G2580_3145_gat), .Y(G3462_3197_gat) );
OR2XL U_g2987 (.A(G7148_3078_ngat), .B(G7147_3142_ngat), .Y(G7149_3198_gat) );
OR2XL U_g2988 (.A(G7060_3079_ngat), .B(G7059_3143_ngat), .Y(G7061_3199_gat) );
AND3XL U_g2989 (.A(G3399_1978_gat), .B(G3417_1979_gat), .C(G2580_3145_gat), .Y(G3464_3200_gat) );
AND2XL U_g2990 (.A(G3417_1979_gat), .B(G2580_3145_gat), .Y(G3465_3201_gat) );
INVXL U_g2991 (.A(G4067_3144_gat), .Y(G4072_3202_gat) );
BUFX20 U_g2992 (.A(G2580_3145_gat), .Y(G4793_3203_gat) );
OR2XL U_g2993 (.A(G6131_3149_ngat), .B(G6128_2611_ngat), .Y(G6133_3204_gat) );
OR2XL U_g2994 (.A(G6073_3150_ngat), .B(G6070_2612_ngat), .Y(G6075_3205_gat) );
OR2XL U_g2995 (.A(G6189_3187_ngat), .B(G6186_2811_ngat), .Y(G6191_3208_gat) );
OR2XL U_g2996 (.A(G6280_3096_ngat), .B(G6279_3155_ngat), .Y(G6281_3209_gat) );
INVXL U_g2997 (.A(G975_3157_gat), .Y(G980_3210_gat) );
INVXL U_g2998 (.A(G4753_3158_gat), .Y(G4759_3211_gat) );
OR2XL U_g2999 (.A(G5542_3102_ngat), .B(G5541_3159_ngat), .Y(G5543_3212_gat) );
OR2XL U_g3000 (.A(G5484_3103_ngat), .B(G5483_3160_ngat), .Y(G5485_3213_gat) );
OR2XL U_g3001 (.A(G2007_3161_gat), .B(G1957_2411_gat), .Y(G2008_3214_gat) );
OR2XL U_g3002 (.A(G5696_2669_ngat), .B(G5689_3164_ngat), .Y(G5698_3215_gat) );
OR2XL U_g3003 (.A(G5608_2670_ngat), .B(G5601_3166_ngat), .Y(G5610_3216_gat) );
OR5XL U_g3004 (.A(G1964_3162_gat), .B(G1962_2086_gat), .C(G1961_2072_gat), .D(G1960_2059_gat), .E(G1880_895_gat), .Y(G4721_3217_gat) );
OR4XL U_g3005 (.A(G1968_3163_gat), .B(G1966_2089_gat), .C(G1965_2074_gat), .D(G1897_900_gat), .Y(G4729_3218_gat) );
INVXL U_g3006 (.A(G5689_3164_gat), .Y(G5695_3219_gat) );
OR3XL U_g3007 (.A(G1971_3165_gat), .B(G1969_2088_gat), .C(G1914_905_gat), .Y(G4737_3220_gat) );
INVXL U_g3008 (.A(G5601_3166_gat), .Y(G5607_3221_gat) );
OR2XL U_g3009 (.A(G1973_3167_gat), .B(G1929_910_gat), .Y(G4745_3222_gat) );
OR2XL U_g3010 (.A(G4720_2430_ngat), .B(G4713_3136_ngat), .Y(G294_3223_gat) );
OR2XL U_g3011 (.A(G4966_1198_ngat), .B(G4959_3170_ngat), .Y(G4968_3224_gat) );
OR2XL U_g3012 (.A(G5007_1201_ngat), .B(G5000_3169_ngat), .Y(G5009_3225_gat) );
INVXL U_g3013 (.A(G5000_3169_gat), .Y(G5006_3226_gat) );
INVXL U_g3014 (.A(G4959_3170_gat), .Y(G4965_3227_gat) );
AND2XL U_g3015 (.A(G955_3172_gat), .B(G933_2683_gat), .Y(G958_3228_gat) );
OR2XL U_g3016 (.A(G1160_3173_gat), .B(G1129_2434_gat), .Y(G1161_3229_gat) );
AND2XL U_g3017 (.A(G3243_3171_gat), .B(G3238_2684_gat), .Y(G3245_3230_gat) );
OR2XL U_g3018 (.A(G5126_2685_ngat), .B(G5119_3175_ngat), .Y(G5128_3231_gat) );
OR2XL U_g3019 (.A(G5038_2686_ngat), .B(G5031_3178_ngat), .Y(G5040_3232_gat) );
OR5XL U_g3020 (.A(G1136_3174_gat), .B(G1134_2131_gat), .C(G1133_2115_gat), .D(G1132_2164_gat), .E(G1050_930_gat), .Y(G4761_3233_gat) );
INVXL U_g3021 (.A(G5119_3175_gat), .Y(G5125_3234_gat) );
OR3XL U_g3022 (.A(G1143_3177_gat), .B(G1141_2133_gat), .C(G1086_935_gat), .Y(G4777_3235_gat) );
INVXL U_g3023 (.A(G5031_3178_gat), .Y(G5037_3236_gat) );
OR2XL U_g3024 (.A(G1145_3179_gat), .B(G1102_940_gat), .Y(G4785_3237_gat) );
OR2XL U_g3025 (.A(G4760_2455_ngat), .B(G4753_3158_ngat), .Y(G323_3238_gat) );
OR2XL U_g3026 (.A(G2866_3115_ngat), .B(G2865_3180_ngat), .Y(G2867_3239_gat) );
OR2XL U_g3027 (.A(G3620_3117_ngat), .B(G3619_3181_ngat), .Y(G3621_3240_gat) );
OR2XL U_g3028 (.A(G3149_3182_ngat), .B(G3136_2475_ngat), .Y(G3150_3241_gat) );
OR4XL U_g3029 (.A(G1140_3176_gat), .B(G1138_2134_gat), .C(G1137_2117_gat), .D(G1068_981_gat), .Y(G4769_3242_gat) );
OR2XL U_g3030 (.A(G4519_3124_ngat), .B(G4518_3183_ngat), .Y(G4520_3243_gat) );
OR2XL U_g3031 (.A(G3617_3126_ngat), .B(G3616_3184_ngat), .Y(G3618_3244_gat) );
OR2XL U_g3032 (.A(G2863_3127_ngat), .B(G2862_3185_ngat), .Y(G2864_3245_gat) );
OR2XL U_g3033 (.A(G4522_3128_ngat), .B(G4521_3186_ngat), .Y(G4523_3246_gat) );
OR2XL U_g3034 (.A(G7002_3138_ngat), .B(G7001_3193_ngat), .Y(G7003_3247_gat) );
OR2XL U_g3035 (.A(G6944_3139_ngat), .B(G6943_3194_ngat), .Y(G6945_3248_gat) );
OR2XL U_g3036 (.A(G3490_3195_gat), .B(G3453_2578_gat), .Y(G3491_3249_gat) );
OR5XL U_g3037 (.A(G3459_3196_gat), .B(G3458_2294_gat), .C(G3457_2282_gat), .D(G3456_2273_gat), .E(G3376_1119_gat), .Y(G4801_3250_gat) );
OR2XL U_g3038 (.A(G7156_2774_ngat), .B(G7149_3198_ngat), .Y(G7158_3251_gat) );
OR2XL U_g3039 (.A(G7068_2775_ngat), .B(G7061_3199_ngat), .Y(G7070_3252_gat) );
OR4XL U_g3040 (.A(G3462_3197_gat), .B(G3461_2297_gat), .C(G3460_2284_gat), .D(G3393_1121_gat), .Y(G4809_3253_gat) );
OR3XL U_g3041 (.A(G3464_3200_gat), .B(G3463_2296_gat), .C(G3410_1123_gat), .Y(G4817_3254_gat) );
INVXL U_g3042 (.A(G7149_3198_gat), .Y(G7155_3255_gat) );
INVXL U_g3043 (.A(G7061_3199_gat), .Y(G7067_3256_gat) );
OR2XL U_g3044 (.A(G3465_3201_gat), .B(G3425_1125_gat), .Y(G4825_3257_gat) );
OR2XL U_g3045 (.A(G4800_2598_ngat), .B(G4793_3203_ngat), .Y(G343_3258_gat) );
INVXL U_g3046 (.A(G4793_3203_gat), .Y(G4799_3259_gat) );
OR2XL U_g3047 (.A(G6134_3146_ngat), .B(G6133_3204_ngat), .Y(G6135_3260_gat) );
OR2XL U_g3048 (.A(G6076_3147_ngat), .B(G6075_3205_ngat), .Y(G6077_3261_gat) );
OR2XL U_g3049 (.A(G6288_2805_ngat), .B(G6281_3209_ngat), .Y(G6290_3262_gat) );
OR2XL U_g3050 (.A(G6192_3154_ngat), .B(G6191_3208_ngat), .Y(G6193_3263_gat) );
INVXL U_g3051 (.A(G6281_3209_gat), .Y(G6287_3264_gat) );
AND4XL U_g3052 (.A(G4523_3246_gat), .B(G4520_3243_gat), .C(G4517_3156_gat), .D(G3615_3168_gat), .Y(G4524_3265_gat) );
AND2XL U_g3053 (.A(G1987_2942_gat), .B(G2008_3214_gat), .Y(G297_3266_gat) );
AND2XL U_g3054 (.A(G1994_2945_gat), .B(G2008_3214_gat), .Y(G300_3267_gat) );
INVXL U_g3055 (.A(G5543_3212_gat), .Y(G5549_3268_gat) );
INVXL U_g3056 (.A(G5485_3213_gat), .Y(G5491_3269_gat) );
AND2XL U_g3057 (.A(G1856_2037_gat), .B(G2008_3214_gat), .Y(G306_3270_gat) );
AND2XL U_g3058 (.A(G2002_2947_gat), .B(G2008_3214_gat), .Y(G303_3271_gat) );
OR2XL U_g3059 (.A(G5550_2401_ngat), .B(G5543_3212_ngat), .Y(G5552_3272_gat) );
OR2XL U_g3060 (.A(G5492_2402_ngat), .B(G5485_3213_ngat), .Y(G5494_3273_gat) );
INVXL U_g3061 (.A(G2008_3214_gat), .Y(G2014_3274_gat) );
OR2XL U_g3062 (.A(G4728_2412_ngat), .B(G4721_3217_ngat), .Y(G309_3275_gat) );
OR2XL U_g3063 (.A(G5695_3219_ngat), .B(G5692_2413_ngat), .Y(G5697_3276_gat) );
OR2XL U_g3064 (.A(G5607_3221_ngat), .B(G5604_2414_ngat), .Y(G5609_3277_gat) );
INVXL U_g3065 (.A(G4721_3217_gat), .Y(G4727_3278_gat) );
OR2XL U_g3066 (.A(G4736_2415_ngat), .B(G4729_3218_ngat), .Y(G312_3279_gat) );
INVXL U_g3067 (.A(G4729_3218_gat), .Y(G4735_3280_gat) );
OR2XL U_g3068 (.A(G4744_2423_ngat), .B(G4737_3220_ngat), .Y(G315_3281_gat) );
INVXL U_g3069 (.A(G4737_3220_gat), .Y(G4743_3282_gat) );
OR2XL U_g3070 (.A(G4752_2425_ngat), .B(G4745_3222_ngat), .Y(G318_3283_gat) );
INVXL U_g3071 (.A(G4745_3222_gat), .Y(G4751_3284_gat) );
OR2XL U_g3072 (.A(G4719_3192_ngat), .B(G4716_2094_ngat), .Y(G293_3285_gat) );
AND2XL U_g3073 (.A(G908_1192_gat), .B(G958_3228_gat), .Y(G275_3286_gat) );
AND2XL U_g3074 (.A(G1161_3229_gat), .B(G1176_1838_gat), .Y(G272_3287_gat) );
OR2XL U_g3075 (.A(G4965_3227_ngat), .B(G4962_919_ngat), .Y(G4967_3288_gat) );
OR2XL U_g3076 (.A(G5006_3226_ngat), .B(G5003_920_ngat), .Y(G5008_3289_gat) );
AND2XL U_g3077 (.A(G1023_1205_gat), .B(G1161_3229_gat), .Y(G1174_3290_gat) );
INVXL U_g3078 (.A(G958_3228_gat), .Y(G961_3291_gat) );
INVXL U_g3079 (.A(G1161_3229_gat), .Y(G1166_3292_gat) );
INVXL U_g3080 (.A(G3245_3230_gat), .Y(G3248_3293_gat) );
OR2XL U_g3081 (.A(G4768_2442_ngat), .B(G4761_3233_ngat), .Y(G326_3294_gat) );
OR2XL U_g3082 (.A(G5125_3234_ngat), .B(G5122_2443_ngat), .Y(G5127_3295_gat) );
OR2XL U_g3083 (.A(G5037_3236_ngat), .B(G5034_2444_ngat), .Y(G5039_3296_gat) );
INVXL U_g3084 (.A(G4761_3233_gat), .Y(G4767_3297_gat) );
OR2XL U_g3085 (.A(G4776_2445_ngat), .B(G4769_3242_ngat), .Y(G329_3298_gat) );
INVXL U_g3086 (.A(G4777_3235_gat), .Y(G4783_3299_gat) );
OR2XL U_g3087 (.A(G4792_2449_ngat), .B(G4785_3237_ngat), .Y(G335_3300_gat) );
INVXL U_g3088 (.A(G4785_3237_gat), .Y(G4791_3301_gat) );
OR2XL U_g3089 (.A(G4759_3211_ngat), .B(G4756_2139_ngat), .Y(G322_3302_gat) );
INVXL U_g3090 (.A(G4769_3242_gat), .Y(G4775_3303_gat) );
OR2XL U_g3091 (.A(G4784_2485_ngat), .B(G4777_3235_ngat), .Y(G332_3304_gat) );
AND2XL U_g3092 (.A(G3150_3241_gat), .B(G3146_2871_gat), .Y(G3152_3305_gat) );
AND2XL U_g3093 (.A(G3223_1698_gat), .B(G3245_3230_gat), .Y(G248_3306_gat) );
AND2XL U_g3094 (.A(G1155_2201_gat), .B(G1161_3229_gat), .Y(G1171_3307_gat) );
AND4XL U_g3095 (.A(G2867_3239_gat), .B(G2864_3245_gat), .C(G2861_3189_gat), .D(G1331_3188_gat), .Y(G2868_3308_gat) );
AND4XL U_g3096 (.A(G3621_3240_gat), .B(G3618_3244_gat), .C(G1334_3190_gat), .D(G1328_3191_gat), .Y(G4443_3309_gat) );
AND2XL U_g3097 (.A(G3248_3293_gat), .B(G3244_1962_gat), .Y(G247_3310_gat) );
AND2XL U_g3098 (.A(G3471_2997_gat), .B(G3491_3249_gat), .Y(G346_3311_gat) );
INVXL U_g3099 (.A(G7003_3247_gat), .Y(G7009_3312_gat) );
INVXL U_g3100 (.A(G6945_3248_gat), .Y(G6951_3313_gat) );
AND2XL U_g3101 (.A(G3478_3001_gat), .B(G3491_3249_gat), .Y(G349_3314_gat) );
OR2XL U_g3102 (.A(G7010_2575_ngat), .B(G7003_3247_ngat), .Y(G7012_3315_gat) );
OR2XL U_g3103 (.A(G6952_2576_ngat), .B(G6945_3248_ngat), .Y(G6954_3316_gat) );
AND2XL U_g3104 (.A(G3350_2261_gat), .B(G3491_3249_gat), .Y(G355_3317_gat) );
AND2XL U_g3105 (.A(G3486_3004_gat), .B(G3491_3249_gat), .Y(G352_3318_gat) );
INVXL U_g3106 (.A(G3491_3249_gat), .Y(G3497_3319_gat) );
OR2XL U_g3107 (.A(G4808_2583_ngat), .B(G4801_3250_ngat), .Y(G358_3320_gat) );
INVXL U_g3108 (.A(G4801_3250_gat), .Y(G4807_3321_gat) );
OR2XL U_g3109 (.A(G7155_3255_ngat), .B(G7152_2584_ngat), .Y(G7157_3322_gat) );
OR2XL U_g3110 (.A(G7067_3256_ngat), .B(G7064_2585_ngat), .Y(G7069_3323_gat) );
OR2XL U_g3111 (.A(G4816_2586_ngat), .B(G4809_3253_ngat), .Y(G361_3324_gat) );
INVXL U_g3112 (.A(G4809_3253_gat), .Y(G4815_3325_gat) );
OR2XL U_g3113 (.A(G4824_2593_ngat), .B(G4817_3254_ngat), .Y(G364_3326_gat) );
INVXL U_g3114 (.A(G4817_3254_gat), .Y(G4823_3327_gat) );
OR2XL U_g3115 (.A(G4832_2597_ngat), .B(G4825_3257_ngat), .Y(G367_3328_gat) );
INVXL U_g3116 (.A(G4825_3257_gat), .Y(G4831_3329_gat) );
OR2XL U_g3117 (.A(G4799_3259_ngat), .B(G4796_2304_ngat), .Y(G342_3330_gat) );
INVXL U_g3118 (.A(G6135_3260_gat), .Y(G6141_3331_gat) );
INVXL U_g3119 (.A(G6077_3261_gat), .Y(G6083_3332_gat) );
OR2XL U_g3120 (.A(G6142_2625_ngat), .B(G6135_3260_ngat), .Y(G6144_3333_gat) );
OR2XL U_g3121 (.A(G6084_2626_ngat), .B(G6077_3261_ngat), .Y(G6086_3334_gat) );
OR2XL U_g3122 (.A(G6287_3264_ngat), .B(G6284_2635_ngat), .Y(G6289_3335_gat) );
OR2XL U_g3123 (.A(G6200_2933_ngat), .B(G6193_3263_ngat), .Y(G6202_3336_gat) );
INVXL U_g3124 (.A(G6193_3263_gat), .Y(G6199_3337_gat) );
AND3XL U_g3125 (.A(G2868_3308_gat), .B(G4524_3265_gat), .C(G4443_3309_gat), .Y(G2881_3339_gat) );
AND2XL U_g3126 (.A(G2014_3274_gat), .B(G1991_3031_gat), .Y(G296_3340_gat) );
AND2XL U_g3127 (.A(G2014_3274_gat), .B(G1998_3036_gat), .Y(G299_3341_gat) );
AND2XL U_g3128 (.A(G2014_3274_gat), .B(G2005_2824_gat), .Y(G302_3342_gat) );
AND2XL U_g3129 (.A(G2014_3274_gat), .B(G1850_1812_gat), .Y(G305_3343_gat) );
OR2XL U_g3130 (.A(G5549_3268_ngat), .B(G5546_2038_ngat), .Y(G5551_3344_gat) );
OR2XL U_g3131 (.A(G5491_3269_ngat), .B(G5488_2039_ngat), .Y(G5493_3345_gat) );
OR2XL U_g3132 (.A(G4727_3278_ngat), .B(G4724_2048_ngat), .Y(G308_3346_gat) );
OR2XL U_g3133 (.A(G5698_3215_ngat), .B(G5697_3276_ngat), .Y(G5699_3347_gat) );
OR2XL U_g3134 (.A(G5610_3216_ngat), .B(G5609_3277_ngat), .Y(G5611_3348_gat) );
OR2XL U_g3135 (.A(G4735_3280_ngat), .B(G4732_2051_ngat), .Y(G311_3349_gat) );
OR2XL U_g3136 (.A(G4743_3282_ngat), .B(G4740_2066_ngat), .Y(G314_3350_gat) );
OR2XL U_g3137 (.A(G4751_3284_ngat), .B(G4748_2075_ngat), .Y(G317_3351_gat) );
AND2XL U_g3138 (.A(G961_3291_gat), .B(G957_1836_gat), .Y(G274_3353_gat) );
AND2XL U_g3139 (.A(G1166_3292_gat), .B(G1117_1193_gat), .Y(G271_3354_gat) );
OR2XL U_g3140 (.A(G4968_3224_ngat), .B(G4967_3288_ngat), .Y(G967_3355_gat) );
OR2XL U_g3141 (.A(G5009_3225_ngat), .B(G5008_3289_ngat), .Y(G971_3356_gat) );
AND2XL U_g3142 (.A(G1166_3292_gat), .B(G1019_923_gat), .Y(G1173_3357_gat) );
OR2XL U_g3143 (.A(G4767_3297_ngat), .B(G4764_2102_ngat), .Y(G325_3358_gat) );
OR2XL U_g3144 (.A(G5128_3231_ngat), .B(G5127_3295_ngat), .Y(G5129_3359_gat) );
OR2XL U_g3145 (.A(G5040_3232_ngat), .B(G5039_3296_ngat), .Y(G5041_3360_gat) );
OR2XL U_g3146 (.A(G4775_3303_ngat), .B(G4772_2105_ngat), .Y(G328_3361_gat) );
OR2XL U_g3147 (.A(G4791_3301_ngat), .B(G4788_2118_ngat), .Y(G334_3362_gat) );
OR2XL U_g3148 (.A(G4783_3299_ngat), .B(G4780_2168_ngat), .Y(G331_3364_gat) );
AND2XL U_g3149 (.A(G3131_2733_gat), .B(G3152_3305_gat), .Y(G251_3365_gat) );
INVXL U_g3150 (.A(G3152_3305_gat), .Y(G3155_3366_gat) );
AND2XL U_g3151 (.A(G1166_3292_gat), .B(G1158_1927_gat), .Y(G1170_3367_gat) );
AND2XL U_g3152 (.A(G3497_3319_gat), .B(G3475_3074_gat), .Y(G345_3370_gat) );
AND2XL U_g3153 (.A(G3497_3319_gat), .B(G3482_3075_gat), .Y(G348_3371_gat) );
AND2XL U_g3154 (.A(G3497_3319_gat), .B(G3489_2906_gat), .Y(G351_3372_gat) );
OR2XL U_g3155 (.A(G7009_3312_ngat), .B(G7006_2259_ngat), .Y(G7011_3373_gat) );
OR2XL U_g3156 (.A(G6951_3313_ngat), .B(G6948_2260_ngat), .Y(G6953_3374_gat) );
AND2XL U_g3157 (.A(G3497_3319_gat), .B(G3344_1970_gat), .Y(G354_3375_gat) );
OR2XL U_g3158 (.A(G4807_3321_ngat), .B(G4804_2266_ngat), .Y(G357_3376_gat) );
OR2XL U_g3159 (.A(G7158_3251_ngat), .B(G7157_3322_ngat), .Y(G7159_3377_gat) );
OR2XL U_g3160 (.A(G7070_3252_ngat), .B(G7069_3323_ngat), .Y(G7071_3378_gat) );
OR2XL U_g3161 (.A(G4815_3325_ngat), .B(G4812_2269_ngat), .Y(G360_3379_gat) );
OR2XL U_g3162 (.A(G4823_3327_ngat), .B(G4820_2281_ngat), .Y(G363_3380_gat) );
OR2XL U_g3163 (.A(G4831_3329_ngat), .B(G4828_2293_ngat), .Y(G366_3381_gat) );
OR2XL U_g3164 (.A(G6141_3331_ngat), .B(G6138_2342_ngat), .Y(G6143_3383_gat) );
OR2XL U_g3165 (.A(G6083_3332_ngat), .B(G6080_2343_ngat), .Y(G6085_3384_gat) );
OR2XL U_g3166 (.A(G6290_3262_ngat), .B(G6289_3335_ngat), .Y(G6291_3385_gat) );
OR2XL U_g3167 (.A(G6199_3337_ngat), .B(G6196_2806_ngat), .Y(G6201_3386_gat) );
OR2XL U_g3168 (.A(G5552_3272_ngat), .B(G5551_3344_ngat), .Y(G5553_3391_gat) );
OR2XL U_g3169 (.A(G5494_3273_ngat), .B(G5493_3345_ngat), .Y(G5495_3392_gat) );
INVXL U_g3170 (.A(G5699_3347_gat), .Y(G5705_3394_gat) );
INVXL U_g3171 (.A(G5611_3348_gat), .Y(G5617_3395_gat) );
OR2XL U_g3172 (.A(G5706_2428_ngat), .B(G5699_3347_ngat), .Y(G5708_3399_gat) );
OR2XL U_g3173 (.A(G5618_2429_ngat), .B(G5611_3348_ngat), .Y(G5620_3400_gat) );
OR2XL U_g3174 (.A(G1174_3290_gat), .B(G1173_3357_gat), .Y(G1175_3403_gat) );
AND3XL U_g3175 (.A(G980_3210_gat), .B(G929_2433_gat), .C(G967_3355_gat), .Y(G992_3404_gat) );
AND3XL U_g3176 (.A(G980_3210_gat), .B(G933_2683_gat), .C(G971_3356_gat), .Y(G991_3405_gat) );
AND3XL U_g3177 (.A(G975_3157_gat), .B(G962_2839_gat), .C(G971_3356_gat), .Y(G993_3406_gat) );
AND3XL U_g3178 (.A(G975_3157_gat), .B(G965_2958_gat), .C(G967_3355_gat), .Y(G994_3407_gat) );
INVXL U_g3179 (.A(G5129_3359_gat), .Y(G5135_3409_gat) );
INVXL U_g3180 (.A(G5041_3360_gat), .Y(G5047_3410_gat) );
OR2XL U_g3181 (.A(G5136_2453_ngat), .B(G5129_3359_ngat), .Y(G5138_3413_gat) );
OR2XL U_g3182 (.A(G5048_2454_ngat), .B(G5041_3360_ngat), .Y(G5050_3414_gat) );
AND3XL U_g3183 (.A(G2881_3339_gat), .B(G2878_386_gat), .C(G2876_389_gat), .Y(G417_3415_gat) );
AND2XL U_g3184 (.A(G3155_3366_gat), .B(G3151_2974_gat), .Y(G250_3417_gat) );
OR2XL U_g3185 (.A(G1171_3307_gat), .B(G1170_3367_gat), .Y(G1172_3419_gat) );
OR2XL U_g3186 (.A(G7012_3315_ngat), .B(G7011_3373_ngat), .Y(G7013_3422_gat) );
OR2XL U_g3187 (.A(G6954_3316_ngat), .B(G6953_3374_ngat), .Y(G6955_3423_gat) );
INVXL U_g3188 (.A(G7159_3377_gat), .Y(G7165_3427_gat) );
INVXL U_g3189 (.A(G7071_3378_gat), .Y(G7077_3428_gat) );
OR2XL U_g3190 (.A(G7166_2599_ngat), .B(G7159_3377_ngat), .Y(G7168_3432_gat) );
OR2XL U_g3191 (.A(G7078_2600_ngat), .B(G7071_3378_ngat), .Y(G7080_3433_gat) );
OR2XL U_g3192 (.A(G6144_3333_ngat), .B(G6143_3383_ngat), .Y(G6145_3434_gat) );
OR2XL U_g3193 (.A(G6086_3334_ngat), .B(G6085_3384_ngat), .Y(G6087_3435_gat) );
INVXL U_g3194 (.A(G6291_3385_gat), .Y(G6297_3436_gat) );
OR2XL U_g3195 (.A(G6202_3336_ngat), .B(G6201_3386_ngat), .Y(G6203_3437_gat) );
OR2XL U_g3196 (.A(G5502_2395_ngat), .B(G5495_3392_ngat), .Y(G5504_3438_gat) );
OR2XL U_g3197 (.A(G5560_2396_ngat), .B(G5553_3391_ngat), .Y(G5562_3439_gat) );
INVXL U_g3198 (.A(G5553_3391_gat), .Y(G5559_3440_gat) );
INVXL U_g3199 (.A(G5495_3392_gat), .Y(G5501_3441_gat) );
OR2XL U_g3200 (.A(G5705_3394_ngat), .B(G5702_2090_ngat), .Y(G5707_3442_gat) );
OR2XL U_g3201 (.A(G5617_3395_ngat), .B(G5614_2091_ngat), .Y(G5619_3443_gat) );
OR4XL U_g3202 (.A(G994_3407_gat), .B(G993_3406_gat), .C(G992_3404_gat), .D(G991_3405_gat), .Y(G5167_3446_gat) );
OR2XL U_g3203 (.A(G5135_3409_ngat), .B(G5132_2135_ngat), .Y(G5137_3447_gat) );
OR2XL U_g3204 (.A(G5047_3410_ngat), .B(G5044_2136_ngat), .Y(G5049_3448_gat) );
OR2XL U_g3205 (.A(G6298_2880_ngat), .B(G6291_3385_ngat), .Y(G6300_3453_gat) );
OR2XL U_g3206 (.A(G6962_2572_ngat), .B(G6955_3423_ngat), .Y(G6964_3454_gat) );
OR2XL U_g3207 (.A(G7020_2573_ngat), .B(G7013_3422_ngat), .Y(G7022_3455_gat) );
INVXL U_g3208 (.A(G7013_3422_gat), .Y(G7019_3456_gat) );
INVXL U_g3209 (.A(G6955_3423_gat), .Y(G6961_3457_gat) );
OR2XL U_g3210 (.A(G7165_3427_ngat), .B(G7162_2305_ngat), .Y(G7167_3458_gat) );
OR2XL U_g3211 (.A(G7077_3428_ngat), .B(G7074_2306_ngat), .Y(G7079_3459_gat) );
OR2XL U_g3212 (.A(G6094_2620_ngat), .B(G6087_3435_ngat), .Y(G6096_3460_gat) );
OR2XL U_g3213 (.A(G6152_2621_ngat), .B(G6145_3434_ngat), .Y(G6154_3461_gat) );
INVXL U_g3214 (.A(G6145_3434_gat), .Y(G6151_3462_gat) );
INVXL U_g3215 (.A(G6087_3435_gat), .Y(G6093_3463_gat) );
INVXL U_g3216 (.A(G6203_3437_gat), .Y(G6209_3464_gat) );
OR2XL U_g3217 (.A(G5501_3441_ngat), .B(G5498_2023_ngat), .Y(G5503_3465_gat) );
OR2XL U_g3218 (.A(G5559_3440_ngat), .B(G5556_2024_ngat), .Y(G5561_3466_gat) );
OR2XL U_g3219 (.A(G5708_3399_ngat), .B(G5707_3442_ngat), .Y(G5709_3467_gat) );
OR2XL U_g3220 (.A(G5620_3400_ngat), .B(G5619_3443_ngat), .Y(G5621_3468_gat) );
INVXL U_g3221 (.A(G5167_3446_gat), .Y(G5173_3469_gat) );
OR2XL U_g3222 (.A(G5138_3413_ngat), .B(G5137_3447_ngat), .Y(G5139_3470_gat) );
OR2XL U_g3223 (.A(G5050_3414_ngat), .B(G5049_3448_ngat), .Y(G5051_3471_gat) );
OR2XL U_g3224 (.A(G6297_3436_ngat), .B(G6294_2746_ngat), .Y(G6299_3472_gat) );
OR2XL U_g3225 (.A(G6210_2881_ngat), .B(G6203_3437_ngat), .Y(G6212_3473_gat) );
OR2XL U_g3226 (.A(G6961_3457_ngat), .B(G6958_2248_ngat), .Y(G6963_3474_gat) );
OR2XL U_g3227 (.A(G7019_3456_ngat), .B(G7016_2249_ngat), .Y(G7021_3475_gat) );
OR2XL U_g3228 (.A(G7168_3432_ngat), .B(G7167_3458_ngat), .Y(G7169_3476_gat) );
OR2XL U_g3229 (.A(G7080_3433_ngat), .B(G7079_3459_ngat), .Y(G7081_3477_gat) );
OR2XL U_g3230 (.A(G6093_3463_ngat), .B(G6090_2328_ngat), .Y(G6095_3478_gat) );
OR2XL U_g3231 (.A(G6151_3462_ngat), .B(G6148_2329_ngat), .Y(G6153_3479_gat) );
OR2XL U_g3232 (.A(G5504_3438_ngat), .B(G5503_3465_ngat), .Y(G5505_3480_gat) );
OR2XL U_g3233 (.A(G5562_3439_ngat), .B(G5561_3466_ngat), .Y(G5563_3481_gat) );
OR2XL U_g3234 (.A(G5628_2426_ngat), .B(G5621_3468_ngat), .Y(G5630_3482_gat) );
OR2XL U_g3235 (.A(G5716_2427_ngat), .B(G5709_3467_ngat), .Y(G5718_3483_gat) );
INVXL U_g3236 (.A(G5709_3467_gat), .Y(G5715_3484_gat) );
INVXL U_g3237 (.A(G5621_3468_gat), .Y(G5627_3485_gat) );
OR2XL U_g3238 (.A(G5058_2451_ngat), .B(G5051_3471_ngat), .Y(G5060_3486_gat) );
OR2XL U_g3239 (.A(G5146_2452_ngat), .B(G5139_3470_ngat), .Y(G5148_3487_gat) );
INVXL U_g3240 (.A(G5139_3470_gat), .Y(G5145_3488_gat) );
INVXL U_g3241 (.A(G5051_3471_gat), .Y(G5057_3489_gat) );
OR2XL U_g3242 (.A(G6300_3453_ngat), .B(G6299_3472_ngat), .Y(G6301_3490_gat) );
OR2XL U_g3243 (.A(G6209_3464_ngat), .B(G6206_2747_ngat), .Y(G6211_3491_gat) );
OR2XL U_g3244 (.A(G6964_3454_ngat), .B(G6963_3474_ngat), .Y(G6965_3492_gat) );
OR2XL U_g3245 (.A(G7022_3455_ngat), .B(G7021_3475_ngat), .Y(G7023_3493_gat) );
OR2XL U_g3246 (.A(G7088_2595_ngat), .B(G7081_3477_ngat), .Y(G7090_3494_gat) );
OR2XL U_g3247 (.A(G7176_2596_ngat), .B(G7169_3476_ngat), .Y(G7178_3495_gat) );
INVXL U_g3248 (.A(G7169_3476_gat), .Y(G7175_3496_gat) );
INVXL U_g3249 (.A(G7081_3477_gat), .Y(G7087_3497_gat) );
OR2XL U_g3250 (.A(G6096_3460_ngat), .B(G6095_3478_ngat), .Y(G6097_3498_gat) );
OR2XL U_g3251 (.A(G6154_3461_ngat), .B(G6153_3479_ngat), .Y(G6155_3499_gat) );
OR2XL U_g3252 (.A(G6308_2647_ngat), .B(G6301_3490_ngat), .Y(G6310_3500_gat) );
OR2XL U_g3253 (.A(G5570_2376_ngat), .B(G5563_3481_ngat), .Y(G5572_3501_gat) );
OR2XL U_g3254 (.A(G5512_2377_ngat), .B(G5505_3480_ngat), .Y(G5514_3502_gat) );
INVXL U_g3255 (.A(G5505_3480_gat), .Y(G5511_3503_gat) );
INVXL U_g3256 (.A(G5563_3481_gat), .Y(G5569_3504_gat) );
OR2XL U_g3257 (.A(G5627_3485_ngat), .B(G5624_2076_ngat), .Y(G5629_3505_gat) );
OR2XL U_g3258 (.A(G5715_3484_ngat), .B(G5712_2077_ngat), .Y(G5717_3506_gat) );
OR2XL U_g3259 (.A(G5057_3489_ngat), .B(G5054_2121_ngat), .Y(G5059_3507_gat) );
OR2XL U_g3260 (.A(G5145_3488_ngat), .B(G5142_2123_ngat), .Y(G5147_3508_gat) );
INVXL U_g3261 (.A(G6301_3490_gat), .Y(G6307_3509_gat) );
OR2XL U_g3262 (.A(G6212_3473_ngat), .B(G6211_3491_ngat), .Y(G6213_3510_gat) );
OR2XL U_g3263 (.A(G7030_2554_ngat), .B(G7023_3493_ngat), .Y(G7032_3511_gat) );
OR2XL U_g3264 (.A(G6972_2555_ngat), .B(G6965_3492_ngat), .Y(G6974_3512_gat) );
INVXL U_g3265 (.A(G6965_3492_gat), .Y(G6971_3513_gat) );
INVXL U_g3266 (.A(G7023_3493_gat), .Y(G7029_3514_gat) );
OR2XL U_g3267 (.A(G7087_3497_ngat), .B(G7084_2290_ngat), .Y(G7089_3515_gat) );
OR2XL U_g3268 (.A(G7175_3496_ngat), .B(G7172_2291_ngat), .Y(G7177_3516_gat) );
OR2XL U_g3269 (.A(G6162_2604_ngat), .B(G6155_3499_ngat), .Y(G6164_3517_gat) );
OR2XL U_g3270 (.A(G6104_2605_ngat), .B(G6097_3498_ngat), .Y(G6106_3518_gat) );
INVXL U_g3271 (.A(G6097_3498_gat), .Y(G6103_3519_gat) );
INVXL U_g3272 (.A(G6155_3499_gat), .Y(G6161_3520_gat) );
OR2XL U_g3273 (.A(G6220_2646_ngat), .B(G6213_3510_ngat), .Y(G6222_3521_gat) );
OR2XL U_g3274 (.A(G6307_3509_ngat), .B(G6304_2370_ngat), .Y(G6309_3522_gat) );
OR2XL U_g3275 (.A(G5569_3504_ngat), .B(G5566_2000_ngat), .Y(G5571_3523_gat) );
OR2XL U_g3276 (.A(G5511_3503_ngat), .B(G5508_2001_ngat), .Y(G5513_3524_gat) );
OR2XL U_g3277 (.A(G5630_3482_ngat), .B(G5629_3505_ngat), .Y(G5631_3525_gat) );
OR2XL U_g3278 (.A(G5718_3483_ngat), .B(G5717_3506_ngat), .Y(G5719_3526_gat) );
OR2XL U_g3279 (.A(G5060_3486_ngat), .B(G5059_3507_ngat), .Y(G5061_3527_gat) );
OR2XL U_g3280 (.A(G5148_3487_ngat), .B(G5147_3508_ngat), .Y(G5149_3528_gat) );
INVXL U_g3281 (.A(G6213_3510_gat), .Y(G6219_3529_gat) );
OR2XL U_g3282 (.A(G7029_3514_ngat), .B(G7026_2225_ngat), .Y(G7031_3530_gat) );
OR2XL U_g3283 (.A(G6971_3513_ngat), .B(G6968_2226_ngat), .Y(G6973_3531_gat) );
OR2XL U_g3284 (.A(G7090_3494_ngat), .B(G7089_3515_ngat), .Y(G7091_3532_gat) );
OR2XL U_g3285 (.A(G7178_3495_ngat), .B(G7177_3516_ngat), .Y(G7179_3533_gat) );
OR2XL U_g3286 (.A(G6161_3520_ngat), .B(G6158_2308_ngat), .Y(G6163_3534_gat) );
OR2XL U_g3287 (.A(G6103_3519_ngat), .B(G6100_2309_ngat), .Y(G6105_3535_gat) );
OR2XL U_g3288 (.A(G6219_3529_ngat), .B(G6216_2369_ngat), .Y(G6221_3536_gat) );
OR2XL U_g3289 (.A(G6310_3500_ngat), .B(G6309_3522_ngat), .Y(G6311_3537_gat) );
OR2XL U_g3290 (.A(G5572_3501_ngat), .B(G5571_3523_ngat), .Y(G5573_3538_gat) );
OR2XL U_g3291 (.A(G5514_3502_ngat), .B(G5513_3524_ngat), .Y(G5515_3539_gat) );
OR2XL U_g3292 (.A(G5726_2408_ngat), .B(G5719_3526_ngat), .Y(G5728_3540_gat) );
OR2XL U_g3293 (.A(G5638_2409_ngat), .B(G5631_3525_ngat), .Y(G5640_3541_gat) );
INVXL U_g3294 (.A(G5631_3525_gat), .Y(G5637_3542_gat) );
INVXL U_g3295 (.A(G5719_3526_gat), .Y(G5725_3543_gat) );
OR2XL U_g3296 (.A(G5156_2439_ngat), .B(G5149_3528_ngat), .Y(G5158_3544_gat) );
OR2XL U_g3297 (.A(G5068_2440_ngat), .B(G5061_3527_ngat), .Y(G5070_3545_gat) );
INVXL U_g3298 (.A(G5061_3527_gat), .Y(G5067_3546_gat) );
INVXL U_g3299 (.A(G5149_3528_gat), .Y(G5155_3547_gat) );
OR2XL U_g3300 (.A(G7032_3511_ngat), .B(G7031_3530_ngat), .Y(G7033_3548_gat) );
OR2XL U_g3301 (.A(G6974_3512_ngat), .B(G6973_3531_ngat), .Y(G6975_3549_gat) );
OR2XL U_g3302 (.A(G7186_2580_ngat), .B(G7179_3533_ngat), .Y(G7188_3550_gat) );
OR2XL U_g3303 (.A(G7098_2581_ngat), .B(G7091_3532_ngat), .Y(G7100_3551_gat) );
INVXL U_g3304 (.A(G7091_3532_gat), .Y(G7097_3552_gat) );
INVXL U_g3305 (.A(G7179_3533_gat), .Y(G7185_3553_gat) );
OR2XL U_g3306 (.A(G6164_3517_ngat), .B(G6163_3534_ngat), .Y(G6165_3554_gat) );
OR2XL U_g3307 (.A(G6106_3518_ngat), .B(G6105_3535_ngat), .Y(G6107_3555_gat) );
OR2XL U_g3308 (.A(G6318_2632_ngat), .B(G6311_3537_ngat), .Y(G6320_3556_gat) );
OR2XL U_g3309 (.A(G6222_3521_ngat), .B(G6221_3536_ngat), .Y(G6223_3557_gat) );
INVXL U_g3310 (.A(G6311_3537_gat), .Y(G6317_3558_gat) );
INVXL U_g3311 (.A(G5573_3538_gat), .Y(G5579_3559_gat) );
INVXL U_g3312 (.A(G5515_3539_gat), .Y(G5521_3560_gat) );
OR2XL U_g3313 (.A(G5522_2389_ngat), .B(G5515_3539_ngat), .Y(G1756_3561_gat) );
OR2XL U_g3314 (.A(G5580_2390_ngat), .B(G5573_3538_ngat), .Y(G1761_3562_gat) );
OR2XL U_g3315 (.A(G5725_3543_ngat), .B(G5722_2044_ngat), .Y(G5727_3563_gat) );
OR2XL U_g3316 (.A(G5637_3542_ngat), .B(G5634_2045_ngat), .Y(G5639_3564_gat) );
OR2XL U_g3317 (.A(G5155_3547_ngat), .B(G5152_2098_ngat), .Y(G5157_3565_gat) );
OR2XL U_g3318 (.A(G5067_3546_ngat), .B(G5064_2099_ngat), .Y(G5069_3566_gat) );
INVXL U_g3319 (.A(G7033_3548_gat), .Y(G7039_3567_gat) );
INVXL U_g3320 (.A(G6975_3549_gat), .Y(G6981_3568_gat) );
OR2XL U_g3321 (.A(G6982_2565_ngat), .B(G6975_3549_ngat), .Y(G4058_3569_gat) );
OR2XL U_g3322 (.A(G7040_2566_ngat), .B(G7033_3548_ngat), .Y(G4063_3570_gat) );
OR2XL U_g3323 (.A(G7185_3553_ngat), .B(G7182_2262_ngat), .Y(G7187_3571_gat) );
OR2XL U_g3324 (.A(G7097_3552_ngat), .B(G7094_2263_ngat), .Y(G7099_3572_gat) );
INVXL U_g3325 (.A(G6165_3554_gat), .Y(G6171_3573_gat) );
INVXL U_g3326 (.A(G6107_3555_gat), .Y(G6113_3574_gat) );
OR2XL U_g3327 (.A(G6114_2615_ngat), .B(G6107_3555_ngat), .Y(G2818_3575_gat) );
OR2XL U_g3328 (.A(G6172_2616_ngat), .B(G6165_3554_ngat), .Y(G2823_3576_gat) );
OR2XL U_g3329 (.A(G6317_3558_ngat), .B(G6314_2346_ngat), .Y(G6319_3577_gat) );
OR2XL U_g3330 (.A(G6230_2633_ngat), .B(G6223_3557_ngat), .Y(G6232_3578_gat) );
INVXL U_g3331 (.A(G6223_3557_gat), .Y(G6229_3579_gat) );
OR2XL U_g3332 (.A(G5521_3560_ngat), .B(G5518_2011_ngat), .Y(G1755_3580_gat) );
OR2XL U_g3333 (.A(G5579_3559_ngat), .B(G5576_2013_ngat), .Y(G1760_3581_gat) );
OR2XL U_g3334 (.A(G5728_3540_ngat), .B(G5727_3563_ngat), .Y(G5729_3582_gat) );
OR2XL U_g3335 (.A(G5640_3541_ngat), .B(G5639_3564_ngat), .Y(G5641_3583_gat) );
OR2XL U_g3336 (.A(G5158_3544_ngat), .B(G5157_3565_ngat), .Y(G5159_3584_gat) );
OR2XL U_g3337 (.A(G5070_3545_ngat), .B(G5069_3566_ngat), .Y(G5071_3585_gat) );
OR2XL U_g3338 (.A(G6981_3568_ngat), .B(G6978_2235_ngat), .Y(G4057_3586_gat) );
OR2XL U_g3339 (.A(G7039_3567_ngat), .B(G7036_2237_ngat), .Y(G4062_3587_gat) );
OR2XL U_g3340 (.A(G7188_3550_ngat), .B(G7187_3571_ngat), .Y(G7189_3588_gat) );
OR2XL U_g3341 (.A(G7100_3551_ngat), .B(G7099_3572_ngat), .Y(G7101_3589_gat) );
OR2XL U_g3342 (.A(G6113_3574_ngat), .B(G6110_2318_ngat), .Y(G2817_3590_gat) );
OR2XL U_g3343 (.A(G6171_3573_ngat), .B(G6168_2320_ngat), .Y(G2822_3591_gat) );
OR2XL U_g3344 (.A(G6320_3556_ngat), .B(G6319_3577_ngat), .Y(G6321_3592_gat) );
OR2XL U_g3345 (.A(G6229_3579_ngat), .B(G6226_2347_ngat), .Y(G6231_3593_gat) );
OR2XL U_g3346 (.A(G1756_3561_ngat), .B(G1755_3580_ngat), .Y(G1757_3594_gat) );
OR2XL U_g3347 (.A(G1761_3562_ngat), .B(G1760_3581_ngat), .Y(G1762_3595_gat) );
INVXL U_g3348 (.A(G5729_3582_gat), .Y(G5735_3596_gat) );
INVXL U_g3349 (.A(G5641_3583_gat), .Y(G5647_3597_gat) );
OR2XL U_g3350 (.A(G5736_2421_ngat), .B(G5729_3582_ngat), .Y(G5660_3598_gat) );
OR2XL U_g3351 (.A(G5648_2422_ngat), .B(G5641_3583_ngat), .Y(G5650_3599_gat) );
INVXL U_g3352 (.A(G5159_3584_gat), .Y(G5165_3600_gat) );
INVXL U_g3353 (.A(G5071_3585_gat), .Y(G5077_3601_gat) );
OR2XL U_g3354 (.A(G5166_2483_ngat), .B(G5159_3584_ngat), .Y(G5090_3602_gat) );
OR2XL U_g3355 (.A(G5078_2484_ngat), .B(G5071_3585_ngat), .Y(G5080_3603_gat) );
OR2XL U_g3356 (.A(G4058_3569_ngat), .B(G4057_3586_ngat), .Y(G4059_3604_gat) );
OR2XL U_g3357 (.A(G4063_3570_ngat), .B(G4062_3587_ngat), .Y(G4064_3605_gat) );
INVXL U_g3358 (.A(G7189_3588_gat), .Y(G7195_3606_gat) );
INVXL U_g3359 (.A(G7101_3589_gat), .Y(G7107_3607_gat) );
OR2XL U_g3360 (.A(G7196_2591_ngat), .B(G7189_3588_ngat), .Y(G7120_3608_gat) );
OR2XL U_g3361 (.A(G7108_2592_ngat), .B(G7101_3589_ngat), .Y(G7110_3609_gat) );
OR2XL U_g3362 (.A(G2818_3575_ngat), .B(G2817_3590_ngat), .Y(G2819_3610_gat) );
OR2XL U_g3363 (.A(G2823_3576_ngat), .B(G2822_3591_ngat), .Y(G2824_3611_gat) );
INVXL U_g3364 (.A(G6321_3592_gat), .Y(G6327_3612_gat) );
OR2XL U_g3365 (.A(G6232_3578_ngat), .B(G6231_3593_ngat), .Y(G6233_3613_gat) );
OR2XL U_g3366 (.A(G6328_2642_ngat), .B(G6321_3592_ngat), .Y(G6252_3614_gat) );
AND3XL U_g3367 (.A(G1771_3137_gat), .B(G1726_2407_gat), .C(G1757_3594_gat), .Y(G1783_3615_gat) );
AND3XL U_g3368 (.A(G1771_3137_gat), .B(G1730_2668_gat), .C(G1762_3595_gat), .Y(G1782_3616_gat) );
AND3XL U_g3369 (.A(G1766_3073_gat), .B(G1751_2828_gat), .C(G1762_3595_gat), .Y(G1784_3617_gat) );
AND3XL U_g3370 (.A(G1766_3073_gat), .B(G1754_2950_gat), .C(G1757_3594_gat), .Y(G1785_3618_gat) );
OR2XL U_g3371 (.A(G5735_3596_ngat), .B(G5732_2063_ngat), .Y(G5659_3619_gat) );
OR2XL U_g3372 (.A(G5647_3597_ngat), .B(G5644_2064_ngat), .Y(G5649_3620_gat) );
OR2XL U_g3373 (.A(G5165_3600_ngat), .B(G5162_2166_ngat), .Y(G5089_3621_gat) );
OR2XL U_g3374 (.A(G5077_3601_ngat), .B(G5074_2167_ngat), .Y(G5079_3622_gat) );
AND3XL U_g3375 (.A(G2828_208_gat), .B(G2813_2930_gat), .C(G2824_3611_gat), .Y(G2846_3623_gat) );
AND3XL U_g3376 (.A(G2828_208_gat), .B(G2816_3019_gat), .C(G2819_3610_gat), .Y(G2847_3624_gat) );
AND3XL U_g3377 (.A(G2833_317_gat), .B(G2784_2802_gat), .C(G2824_3611_gat), .Y(G2844_3625_gat) );
AND3XL U_g3378 (.A(G2833_317_gat), .B(G2780_2629_gat), .C(G2819_3610_gat), .Y(G2845_3626_gat) );
AND3XL U_g3379 (.A(G4072_3202_gat), .B(G4028_2579_gat), .C(G4059_3604_gat), .Y(G4084_3627_gat) );
AND3XL U_g3380 (.A(G4072_3202_gat), .B(G4032_2773_gat), .C(G4064_3605_gat), .Y(G4083_3628_gat) );
AND3XL U_g3381 (.A(G4067_3144_gat), .B(G4053_2910_gat), .C(G4064_3605_gat), .Y(G4085_3629_gat) );
AND3XL U_g3382 (.A(G4067_3144_gat), .B(G4056_3005_gat), .C(G4059_3604_gat), .Y(G4086_3630_gat) );
OR2XL U_g3383 (.A(G7195_3606_ngat), .B(G7192_2278_ngat), .Y(G7119_3631_gat) );
OR2XL U_g3384 (.A(G7107_3607_ngat), .B(G7104_2279_ngat), .Y(G7109_3632_gat) );
INVXL U_g3385 (.A(G6233_3613_gat), .Y(G6239_3633_gat) );
OR2XL U_g3386 (.A(G6327_3612_ngat), .B(G6324_2359_ngat), .Y(G6251_3634_gat) );
OR2XL U_g3387 (.A(G6240_2643_ngat), .B(G6233_3613_ngat), .Y(G6242_3635_gat) );
OR4XL U_g3388 (.A(G1785_3618_gat), .B(G1784_3617_gat), .C(G1783_3615_gat), .D(G1782_3616_gat), .Y(G5737_3636_gat) );
OR2XL U_g3389 (.A(G5660_3598_ngat), .B(G5659_3619_ngat), .Y(G5661_3637_gat) );
OR2XL U_g3390 (.A(G5650_3599_ngat), .B(G5649_3620_ngat), .Y(G5651_3638_gat) );
OR2XL U_g3391 (.A(G5090_3602_ngat), .B(G5089_3621_ngat), .Y(G5091_3639_gat) );
OR2XL U_g3392 (.A(G5080_3603_ngat), .B(G5079_3622_ngat), .Y(G5081_3640_gat) );
OR4XL U_g3393 (.A(G2847_3624_gat), .B(G2846_3623_gat), .C(G2845_3626_gat), .D(G2844_3625_gat), .Y(G6329_3641_gat) );
OR4XL U_g3394 (.A(G4086_3630_gat), .B(G4085_3629_gat), .C(G4084_3627_gat), .D(G4083_3628_gat), .Y(G7197_3642_gat) );
OR2XL U_g3395 (.A(G7120_3608_ngat), .B(G7119_3631_ngat), .Y(G7121_3643_gat) );
OR2XL U_g3396 (.A(G7110_3609_ngat), .B(G7109_3632_ngat), .Y(G7111_3644_gat) );
OR2XL U_g3397 (.A(G6252_3614_ngat), .B(G6251_3634_ngat), .Y(G6253_3645_gat) );
OR2XL U_g3398 (.A(G6239_3633_ngat), .B(G6236_2360_ngat), .Y(G6241_3646_gat) );
INVXL U_g3399 (.A(G5737_3636_gat), .Y(G5743_3647_gat) );
OR2XL U_g3400 (.A(G5668_2416_ngat), .B(G5661_3637_ngat), .Y(G1779_3648_gat) );
OR2XL U_g3401 (.A(G5658_2417_ngat), .B(G5651_3638_ngat), .Y(G1776_3649_gat) );
INVXL U_g3402 (.A(G5661_3637_gat), .Y(G5667_3650_gat) );
INVXL U_g3403 (.A(G5651_3638_gat), .Y(G5657_3651_gat) );
OR2XL U_g3404 (.A(G5098_2446_ngat), .B(G5091_3639_ngat), .Y(G988_3652_gat) );
OR2XL U_g3405 (.A(G5088_2447_ngat), .B(G5081_3640_ngat), .Y(G985_3653_gat) );
INVXL U_g3406 (.A(G5091_3639_gat), .Y(G5097_3654_gat) );
INVXL U_g3407 (.A(G5081_3640_gat), .Y(G5087_3655_gat) );
INVXL U_g3408 (.A(G6329_3641_gat), .Y(G6335_3656_gat) );
INVXL U_g3409 (.A(G7197_3642_gat), .Y(G7203_3657_gat) );
OR2XL U_g3410 (.A(G7128_2587_ngat), .B(G7121_3643_ngat), .Y(G4080_3658_gat) );
OR2XL U_g3411 (.A(G7118_2588_ngat), .B(G7111_3644_ngat), .Y(G4077_3659_gat) );
INVXL U_g3412 (.A(G7121_3643_gat), .Y(G7127_3660_gat) );
INVXL U_g3413 (.A(G7111_3644_gat), .Y(G7117_3661_gat) );
OR2XL U_g3414 (.A(G6260_2636_ngat), .B(G6253_3645_ngat), .Y(G2841_3662_gat) );
INVXL U_g3415 (.A(G6253_3645_gat), .Y(G6259_3663_gat) );
OR2XL U_g3416 (.A(G6242_3635_ngat), .B(G6241_3646_ngat), .Y(G6243_3664_gat) );
OR2XL U_g3417 (.A(G5667_3650_ngat), .B(G5664_2052_ngat), .Y(G1778_3665_gat) );
OR2XL U_g3418 (.A(G5657_3651_ngat), .B(G5654_2054_ngat), .Y(G1775_3666_gat) );
OR2XL U_g3419 (.A(G5097_3654_ngat), .B(G5094_2106_ngat), .Y(G987_3667_gat) );
OR2XL U_g3420 (.A(G5087_3655_ngat), .B(G5084_2108_ngat), .Y(G984_3668_gat) );
OR2XL U_g3421 (.A(G7127_3660_ngat), .B(G7124_2270_ngat), .Y(G4079_3669_gat) );
OR2XL U_g3422 (.A(G7117_3661_ngat), .B(G7114_2272_ngat), .Y(G4076_3670_gat) );
OR2XL U_g3423 (.A(G6259_3663_ngat), .B(G6256_2350_ngat), .Y(G2840_3671_gat) );
OR2XL U_g3424 (.A(G6250_2638_ngat), .B(G6243_3664_ngat), .Y(G2838_3672_gat) );
INVXL U_g3425 (.A(G6243_3664_gat), .Y(G6249_3673_gat) );
OR2XL U_g3426 (.A(G1779_3648_ngat), .B(G1778_3665_ngat), .Y(G1780_3674_gat) );
OR2XL U_g3427 (.A(G1776_3649_ngat), .B(G1775_3666_ngat), .Y(G1777_3675_gat) );
OR2XL U_g3428 (.A(G988_3652_ngat), .B(G987_3667_ngat), .Y(G989_3676_gat) );
OR2XL U_g3429 (.A(G985_3653_ngat), .B(G984_3668_ngat), .Y(G986_3677_gat) );
AND2XL U_g3430 (.A(G1777_3675_gat), .B(G1766_3073_gat), .Y(G1787_3678_gat) );
OR2XL U_g3431 (.A(G4080_3658_ngat), .B(G4079_3669_ngat), .Y(G4081_3679_gat) );
OR2XL U_g3432 (.A(G4077_3659_ngat), .B(G4076_3670_ngat), .Y(G4078_3680_gat) );
OR2XL U_g3433 (.A(G2841_3662_ngat), .B(G2840_3671_ngat), .Y(G2842_3681_gat) );
OR2XL U_g3434 (.A(G6249_3673_ngat), .B(G6246_2351_ngat), .Y(G2837_3682_gat) );
AND2XL U_g3435 (.A(G986_3677_gat), .B(G975_3157_gat), .Y(G996_3683_gat) );
INVXL U_g3436 (.A(G1780_3674_gat), .Y(G1781_3684_gat) );
INVXL U_g3437 (.A(G989_3676_gat), .Y(G990_3685_gat) );
AND2XL U_g3438 (.A(G1771_3137_gat), .B(G1781_3684_gat), .Y(G1786_3686_gat) );
INVXL U_g3439 (.A(G4081_3679_gat), .Y(G4082_3687_gat) );
AND2XL U_g3440 (.A(G4078_3680_gat), .B(G4067_3144_gat), .Y(G4088_3688_gat) );
INVXL U_g3441 (.A(G2842_3681_gat), .Y(G2843_3689_gat) );
OR2XL U_g3442 (.A(G2838_3672_ngat), .B(G2837_3682_ngat), .Y(G2839_3690_gat) );
AND2XL U_g3443 (.A(G980_3210_gat), .B(G990_3685_gat), .Y(G995_3691_gat) );
AND2XL U_g3444 (.A(G2839_3690_gat), .B(G2828_208_gat), .Y(G2849_3692_gat) );
AND2XL U_g3445 (.A(G2833_317_gat), .B(G2843_3689_gat), .Y(G2848_3693_gat) );
OR2XL U_g3446 (.A(G1787_3678_gat), .B(G1786_3686_gat), .Y(G5740_3694_gat) );
AND2XL U_g3447 (.A(G4072_3202_gat), .B(G4082_3687_gat), .Y(G4087_3695_gat) );
OR2XL U_g3448 (.A(G996_3683_gat), .B(G995_3691_gat), .Y(G5170_3696_gat) );
OR2XL U_g3449 (.A(G2849_3692_gat), .B(G2848_3693_gat), .Y(G6332_3697_gat) );
INVXL U_g3450 (.A(G5740_3694_gat), .Y(G5744_3698_gat) );
OR2XL U_g3451 (.A(G4088_3688_gat), .B(G4087_3695_gat), .Y(G7200_3699_gat) );
INVXL U_g3452 (.A(G5170_3696_gat), .Y(G5174_3700_gat) );
OR2XL U_g3453 (.A(G5743_3647_ngat), .B(G5740_3694_ngat), .Y(G1791_3701_gat) );
OR2XL U_g3454 (.A(G5173_3469_ngat), .B(G5170_3696_ngat), .Y(G1003_3702_gat) );
OR2XL U_g3455 (.A(G6335_3656_ngat), .B(G6332_3697_ngat), .Y(G2855_3703_gat) );
INVXL U_g3456 (.A(G6332_3697_gat), .Y(G6336_3704_gat) );
OR2XL U_g3457 (.A(G7203_3657_ngat), .B(G7200_3699_ngat), .Y(G4092_3705_gat) );
INVXL U_g3458 (.A(G7200_3699_gat), .Y(G7204_3706_gat) );
OR2XL U_g3459 (.A(G5744_3698_ngat), .B(G5737_3636_ngat), .Y(G1792_3707_gat) );
OR2XL U_g3460 (.A(G5174_3700_ngat), .B(G5167_3446_ngat), .Y(G1004_3708_gat) );
OR2XL U_g3461 (.A(G6336_3704_ngat), .B(G6329_3641_ngat), .Y(G2856_3709_gat) );
OR2XL U_g3462 (.A(G7204_3706_ngat), .B(G7197_3642_ngat), .Y(G4093_3710_gat) );
OR2XL U_g3463 (.A(G1792_3707_ngat), .B(G1791_3701_ngat), .Y(G320_3711_gat) );
OR2XL U_g3464 (.A(G1004_3708_ngat), .B(G1003_3702_ngat), .Y(G337_3712_gat) );
OR2XL U_g3465 (.A(G2856_3709_ngat), .B(G2855_3703_ngat), .Y(G398_3713_gat) );
OR2XL U_g3466 (.A(G4093_3710_ngat), .B(G4092_3705_ngat), .Y(G369_3714_gat) );
BUFX20 U_g3467 (.A(GIN_339_164_gat), .Y(G339_164_gat) );
BUFX20 U_g3468 (.A(G1_0_gat), .Y(G2_313_gat) );
BUFX20 U_g3469 (.A(G1_0_gat), .Y(G3_312_gat) );
BUFX20 U_g3470 (.A(G1459_167_gat), .Y(G450_288_gat) );
BUFX20 U_g3471 (.A(G1469_169_gat), .Y(G448_284_gat) );
BUFX20 U_g3472 (.A(G1480_170_gat), .Y(G444_282_gat) );
BUFX20 U_g3473 (.A(G1486_171_gat), .Y(G442_280_gat) );
BUFX20 U_g3474 (.A(G1492_172_gat), .Y(G440_277_gat) );
BUFX20 U_g3475 (.A(G1496_173_gat), .Y(G438_274_gat) );
BUFX20 U_g3476 (.A(G2208_175_gat), .Y(G496_271_gat) );
BUFX20 U_g3477 (.A(G2218_177_gat), .Y(G494_267_gat) );
BUFX20 U_g3478 (.A(G2224_178_gat), .Y(G492_265_gat) );
BUFX20 U_g3479 (.A(G2230_179_gat), .Y(G490_263_gat) );
BUFX20 U_g3480 (.A(G2236_180_gat), .Y(G488_260_gat) );
BUFX20 U_g3481 (.A(G2239_181_gat), .Y(G486_258_gat) );
BUFX20 U_g3482 (.A(G2247_182_gat), .Y(G484_256_gat) );
BUFX20 U_g3483 (.A(G2253_183_gat), .Y(G482_253_gat) );
BUFX20 U_g3484 (.A(G2256_184_gat), .Y(G480_250_gat) );
BUFX20 U_g3485 (.A(G3698_185_gat), .Y(G560_248_gat) );
BUFX20 U_g3486 (.A(G3701_186_gat), .Y(G542_246_gat) );
BUFX20 U_g3487 (.A(G3705_187_gat), .Y(G558_244_gat) );
BUFX20 U_g3488 (.A(G3711_188_gat), .Y(G556_242_gat) );
BUFX20 U_g3489 (.A(G3717_189_gat), .Y(G554_240_gat) );
BUFX20 U_g3490 (.A(G3723_190_gat), .Y(G552_238_gat) );
BUFX20 U_g3491 (.A(G3729_191_gat), .Y(G550_236_gat) );
BUFX20 U_g3492 (.A(G3737_192_gat), .Y(G548_234_gat) );
BUFX20 U_g3493 (.A(G3743_193_gat), .Y(G546_232_gat) );
BUFX20 U_g3494 (.A(G3749_194_gat), .Y(G544_230_gat) );
BUFX20 U_g3495 (.A(G4393_195_gat), .Y(G540_227_gat) );
BUFX20 U_g3496 (.A(G4400_197_gat), .Y(G538_224_gat) );
BUFX20 U_g3497 (.A(G4405_198_gat), .Y(G536_222_gat) );
BUFX20 U_g3498 (.A(G4410_199_gat), .Y(G534_220_gat) );
BUFX20 U_g3499 (.A(G4415_200_gat), .Y(G532_218_gat) );
BUFX20 U_g3500 (.A(G4420_201_gat), .Y(G530_216_gat) );
BUFX20 U_g3501 (.A(G4427_202_gat), .Y(G528_214_gat) );
BUFX20 U_g3502 (.A(G4432_203_gat), .Y(G526_212_gat) );
BUFX20 U_g3503 (.A(G4437_204_gat), .Y(G524_210_gat) );
BUFX20 U_g3504 (.A(G1462_168_gat), .Y(G436_286_gat) );
BUFX20 U_g3505 (.A(G2211_176_gat), .Y(G478_269_gat) );
BUFX20 U_g3506 (.A(G4394_196_gat), .Y(G522_226_gat) );
BUFX20 U_g3507 (.A(G1172_3419_gat), .Y(G422_3451_gat) );
BUFX20 U_g3508 (.A(G1172_3419_gat), .Y(G469_3452_gat) );
BUFX20 U_g3509 (.A(G1175_3403_gat), .Y(G419_3444_gat) );
BUFX20 U_g3510 (.A(G1175_3403_gat), .Y(G471_3445_gat) );
INVXL U_g3511 (.A(G400_297_gat), .Y(G400_297_ngat) );
INVXL U_g3512 (.A(G401_310_gat), .Y(G401_310_ngat) );
INVXL U_g3513 (.A(G1197_165_gat), .Y(G1197_165_ngat) );
INVXL U_g3514 (.A(G574_308_gat), .Y(G574_308_ngat) );
INVXL U_g3515 (.A(G1184_294_gat), .Y(G1184_294_ngat) );
INVXL U_g3516 (.A(G575_309_gat), .Y(G575_309_ngat) );
INVXL U_g3517 (.A(G371_2754_gat), .Y(G371_2754_ngat) );
INVXL U_g3518 (.A(G372_2890_gat), .Y(G372_2890_ngat) );
INVXL U_g3519 (.A(G386_3020_gat), .Y(G386_3020_ngat) );
INVXL U_g3520 (.A(G387_2931_gat), .Y(G387_2931_ngat) );
INVXL U_g3521 (.A(G389_3021_gat), .Y(G389_3021_ngat) );
INVXL U_g3522 (.A(G390_2934_gat), .Y(G390_2934_ngat) );
INVXL U_g3523 (.A(G392_3022_gat), .Y(G392_3022_ngat) );
INVXL U_g3524 (.A(G393_2937_gat), .Y(G393_2937_ngat) );
INVXL U_g3525 (.A(G395_3023_gat), .Y(G395_3023_ngat) );
INVXL U_g3526 (.A(G396_2941_gat), .Y(G396_2941_ngat) );
INVXL U_g3527 (.A(G293_3285_gat), .Y(G293_3285_ngat) );
INVXL U_g3528 (.A(G294_3223_gat), .Y(G294_3223_ngat) );
INVXL U_g3529 (.A(G322_3302_gat), .Y(G322_3302_ngat) );
INVXL U_g3530 (.A(G323_3238_gat), .Y(G323_3238_ngat) );
INVXL U_g3531 (.A(G308_3346_gat), .Y(G308_3346_ngat) );
INVXL U_g3532 (.A(G309_3275_gat), .Y(G309_3275_ngat) );
INVXL U_g3533 (.A(G311_3349_gat), .Y(G311_3349_ngat) );
INVXL U_g3534 (.A(G312_3279_gat), .Y(G312_3279_ngat) );
INVXL U_g3535 (.A(G314_3350_gat), .Y(G314_3350_ngat) );
INVXL U_g3536 (.A(G315_3281_gat), .Y(G315_3281_ngat) );
INVXL U_g3537 (.A(G317_3351_gat), .Y(G317_3351_ngat) );
INVXL U_g3538 (.A(G318_3283_gat), .Y(G318_3283_ngat) );
INVXL U_g3539 (.A(G325_3358_gat), .Y(G325_3358_ngat) );
INVXL U_g3540 (.A(G326_3294_gat), .Y(G326_3294_ngat) );
INVXL U_g3541 (.A(G328_3361_gat), .Y(G328_3361_ngat) );
INVXL U_g3542 (.A(G329_3298_gat), .Y(G329_3298_ngat) );
INVXL U_g3543 (.A(G331_3364_gat), .Y(G331_3364_ngat) );
INVXL U_g3544 (.A(G332_3304_gat), .Y(G332_3304_ngat) );
INVXL U_g3545 (.A(G334_3362_gat), .Y(G334_3362_ngat) );
INVXL U_g3546 (.A(G335_3300_gat), .Y(G335_3300_ngat) );
INVXL U_g3547 (.A(G342_3330_gat), .Y(G342_3330_ngat) );
INVXL U_g3548 (.A(G343_3258_gat), .Y(G343_3258_ngat) );
INVXL U_g3549 (.A(G357_3376_gat), .Y(G357_3376_ngat) );
INVXL U_g3550 (.A(G358_3320_gat), .Y(G358_3320_ngat) );
INVXL U_g3551 (.A(G360_3379_gat), .Y(G360_3379_ngat) );
INVXL U_g3552 (.A(G361_3324_gat), .Y(G361_3324_ngat) );
INVXL U_g3553 (.A(G363_3380_gat), .Y(G363_3380_ngat) );
INVXL U_g3554 (.A(G364_3326_gat), .Y(G364_3326_ngat) );
INVXL U_g3555 (.A(G366_3381_gat), .Y(G366_3381_ngat) );
INVXL U_g3556 (.A(G367_3328_gat), .Y(G367_3328_ngat) );
INVXL U_g3557 (.A(G4528_206_gat), .Y(G4528_206_ngat) );
INVXL U_g3558 (.A(G1496_173_gat), .Y(G1496_173_ngat) );
INVXL U_g3559 (.A(G12_3_gat), .Y(G12_3_ngat) );
INVXL U_g3560 (.A(G9_2_gat), .Y(G9_2_ngat) );
INVXL U_g3561 (.A(G2207_272_gat), .Y(G2207_272_ngat) );
INVXL U_g3562 (.A(G1198_299_gat), .Y(G1198_299_ngat) );
INVXL U_g3563 (.A(G1519_374_gat), .Y(G1519_374_ngat) );
INVXL U_g3564 (.A(G6511_429_gat), .Y(G6511_429_ngat) );
INVXL U_g3565 (.A(G6518_558_gat), .Y(G6518_558_ngat) );
INVXL U_g3566 (.A(G5175_372_gat), .Y(G5175_372_ngat) );
INVXL U_g3567 (.A(G5182_563_gat), .Y(G5182_563_ngat) );
INVXL U_g3568 (.A(G4873_373_gat), .Y(G4873_373_ngat) );
INVXL U_g3569 (.A(G4880_566_gat), .Y(G4880_566_ngat) );
INVXL U_g3570 (.A(G4913_497_gat), .Y(G4913_497_ngat) );
INVXL U_g3571 (.A(G4920_565_gat), .Y(G4920_565_ngat) );
INVXL U_g3572 (.A(G5183_498_gat), .Y(G5183_498_ngat) );
INVXL U_g3573 (.A(G5190_562_gat), .Y(G5190_562_ngat) );
INVXL U_g3574 (.A(G5178_399_gat), .Y(G5178_399_ngat) );
INVXL U_g3575 (.A(G5181_494_gat), .Y(G5181_494_ngat) );
INVXL U_g3576 (.A(G4876_401_gat), .Y(G4876_401_ngat) );
INVXL U_g3577 (.A(G4879_495_gat), .Y(G4879_495_ngat) );
INVXL U_g3578 (.A(G1005_721_gat), .Y(G1005_721_ngat) );
INVXL U_g3579 (.A(G1006_602_gat), .Y(G1006_602_ngat) );
INVXL U_g3580 (.A(G763_723_gat), .Y(G763_723_ngat) );
INVXL U_g3581 (.A(G764_603_gat), .Y(G764_603_ngat) );
INVXL U_g3582 (.A(G6551_599_gat), .Y(G6551_599_ngat) );
INVXL U_g3583 (.A(G6558_556_gat), .Y(G6558_556_ngat) );
INVXL U_g3584 (.A(G6514_397_gat), .Y(G6514_397_ngat) );
INVXL U_g3585 (.A(G6517_598_gat), .Y(G6517_598_ngat) );
INVXL U_g3586 (.A(G5186_398_gat), .Y(G5186_398_ngat) );
INVXL U_g3587 (.A(G5189_607_gat), .Y(G5189_607_ngat) );
INVXL U_g3588 (.A(G4916_400_gat), .Y(G4916_400_ngat) );
INVXL U_g3589 (.A(G4919_605_gat), .Y(G4919_605_ngat) );
INVXL U_g3590 (.A(G3168_828_gat), .Y(G3168_828_ngat) );
INVXL U_g3591 (.A(G3169_597_gat), .Y(G3169_597_ngat) );
INVXL U_g3592 (.A(G737_854_gat), .Y(G737_854_ngat) );
INVXL U_g3593 (.A(G2241_257_gat), .Y(G2241_257_ngat) );
INVXL U_g3594 (.A(G2213_268_gat), .Y(G2213_268_ngat) );
INVXL U_g3595 (.A(G1399_820_gat), .Y(G1399_820_ngat) );
INVXL U_g3596 (.A(G885_832_gat), .Y(G885_832_ngat) );
INVXL U_g3597 (.A(G886_604_gat), .Y(G886_604_ngat) );
INVXL U_g3598 (.A(G1017_831_gat), .Y(G1017_831_ngat) );
INVXL U_g3599 (.A(G1018_606_gat), .Y(G1018_606_ngat) );
INVXL U_g3600 (.A(G1464_285_gat), .Y(G1464_285_ngat) );
INVXL U_g3601 (.A(G2933_861_gat), .Y(G2933_861_ngat) );
INVXL U_g3602 (.A(G6554_396_gat), .Y(G6554_396_ngat) );
INVXL U_g3603 (.A(G6557_741_gat), .Y(G6557_741_ngat) );
INVXL U_g3604 (.A(G4422_215_gat), .Y(G4422_215_ngat) );
INVXL U_g3605 (.A(G3821_1034_gat), .Y(G3821_1034_ngat) );
INVXL U_g3606 (.A(G4396_225_gat), .Y(G4396_225_ngat) );
INVXL U_g3607 (.A(G2179_977_gat), .Y(G2179_977_ngat) );
INVXL U_g3608 (.A(G3731_235_gat), .Y(G3731_235_ngat) );
INVXL U_g3609 (.A(G2091_969_gat), .Y(G2091_969_ngat) );
INVXL U_g3610 (.A(G5396_1084_gat), .Y(G5396_1084_ngat) );
INVXL U_g3611 (.A(G5399_466_gat), .Y(G5399_466_ngat) );
INVXL U_g3612 (.A(G5748_1085_gat), .Y(G5748_1085_ngat) );
INVXL U_g3613 (.A(G5751_467_gat), .Y(G5751_467_ngat) );
INVXL U_g3614 (.A(G5756_1086_gat), .Y(G5756_1086_ngat) );
INVXL U_g3615 (.A(G5759_469_gat), .Y(G5759_469_ngat) );
INVXL U_g3616 (.A(G5404_1087_gat), .Y(G5404_1087_ngat) );
INVXL U_g3617 (.A(G5407_470_gat), .Y(G5407_470_ngat) );
INVXL U_g3618 (.A(G5412_1076_gat), .Y(G5412_1076_ngat) );
INVXL U_g3619 (.A(G5415_472_gat), .Y(G5415_472_ngat) );
INVXL U_g3620 (.A(G5764_1075_gat), .Y(G5764_1075_ngat) );
INVXL U_g3621 (.A(G5767_473_gat), .Y(G5767_473_ngat) );
INVXL U_g3622 (.A(G5772_1078_gat), .Y(G5772_1078_ngat) );
INVXL U_g3623 (.A(G5775_474_gat), .Y(G5775_474_ngat) );
INVXL U_g3624 (.A(G5452_1077_gat), .Y(G5452_1077_ngat) );
INVXL U_g3625 (.A(G5455_475_gat), .Y(G5455_475_ngat) );
INVXL U_g3626 (.A(G5420_1082_gat), .Y(G5420_1082_ngat) );
INVXL U_g3627 (.A(G5423_478_gat), .Y(G5423_478_ngat) );
INVXL U_g3628 (.A(G5780_1081_gat), .Y(G5780_1081_ngat) );
INVXL U_g3629 (.A(G5783_479_gat), .Y(G5783_479_ngat) );
INVXL U_g3630 (.A(G5788_964_gat), .Y(G5788_964_ngat) );
INVXL U_g3631 (.A(G5791_480_gat), .Y(G5791_480_ngat) );
INVXL U_g3632 (.A(G5428_963_gat), .Y(G5428_963_ngat) );
INVXL U_g3633 (.A(G5431_481_gat), .Y(G5431_481_ngat) );
INVXL U_g3634 (.A(G5436_961_gat), .Y(G5436_961_ngat) );
INVXL U_g3635 (.A(G5439_484_gat), .Y(G5439_484_ngat) );
INVXL U_g3636 (.A(G5796_960_gat), .Y(G5796_960_ngat) );
INVXL U_g3637 (.A(G5799_485_gat), .Y(G5799_485_ngat) );
INVXL U_g3638 (.A(G5804_958_gat), .Y(G5804_958_ngat) );
INVXL U_g3639 (.A(G5807_486_gat), .Y(G5807_486_ngat) );
INVXL U_g3640 (.A(G5444_957_gat), .Y(G5444_957_ngat) );
INVXL U_g3641 (.A(G5447_487_gat), .Y(G5447_487_ngat) );
INVXL U_g3642 (.A(G5460_967_gat), .Y(G5460_967_ngat) );
INVXL U_g3643 (.A(G5463_489_gat), .Y(G5463_489_ngat) );
INVXL U_g3644 (.A(G7463_913_gat), .Y(G7463_913_ngat) );
INVXL U_g3645 (.A(G7470_915_gat), .Y(G7470_915_ngat) );
INVXL U_g3646 (.A(G5812_966_gat), .Y(G5812_966_ngat) );
INVXL U_g3647 (.A(G5815_491_gat), .Y(G5815_491_ngat) );
INVXL U_g3648 (.A(G6711_772_gat), .Y(G6711_772_ngat) );
INVXL U_g3649 (.A(G6718_921_gat), .Y(G6718_921_ngat) );
INVXL U_g3650 (.A(G777_370_gat), .Y(G777_370_ngat) );
INVXL U_g3651 (.A(G915_1029_gat), .Y(G915_1029_ngat) );
INVXL U_g3652 (.A(G6714_775_gat), .Y(G6714_775_ngat) );
INVXL U_g3653 (.A(G6717_916_gat), .Y(G6717_916_ngat) );
INVXL U_g3654 (.A(G4884_1105_gat), .Y(G4884_1105_ngat) );
INVXL U_g3655 (.A(G4887_500_gat), .Y(G4887_500_ngat) );
INVXL U_g3656 (.A(G5194_1106_gat), .Y(G5194_1106_ngat) );
INVXL U_g3657 (.A(G5197_501_gat), .Y(G5197_501_ngat) );
INVXL U_g3658 (.A(G5202_1089_gat), .Y(G5202_1089_ngat) );
INVXL U_g3659 (.A(G5205_502_gat), .Y(G5205_502_ngat) );
INVXL U_g3660 (.A(G4892_1090_gat), .Y(G4892_1090_ngat) );
INVXL U_g3661 (.A(G4895_503_gat), .Y(G4895_503_ngat) );
INVXL U_g3662 (.A(G5218_1095_gat), .Y(G5218_1095_ngat) );
INVXL U_g3663 (.A(G5221_505_gat), .Y(G5221_505_ngat) );
INVXL U_g3664 (.A(G4908_1096_gat), .Y(G4908_1096_ngat) );
INVXL U_g3665 (.A(G4911_507_gat), .Y(G4911_507_ngat) );
INVXL U_g3666 (.A(G4924_1099_gat), .Y(G4924_1099_ngat) );
INVXL U_g3667 (.A(G4927_508_gat), .Y(G4927_508_ngat) );
INVXL U_g3668 (.A(G6687_943_gat), .Y(G6687_943_ngat) );
INVXL U_g3669 (.A(G6694_945_gat), .Y(G6694_945_ngat) );
INVXL U_g3670 (.A(G5226_1100_gat), .Y(G5226_1100_ngat) );
INVXL U_g3671 (.A(G5229_510_gat), .Y(G5229_510_ngat) );
INVXL U_g3672 (.A(G7293_953_gat), .Y(G7293_953_ngat) );
INVXL U_g3673 (.A(G7300_946_gat), .Y(G7300_946_ngat) );
INVXL U_g3674 (.A(G5315_965_gat), .Y(G5315_965_ngat) );
INVXL U_g3675 (.A(G5322_955_gat), .Y(G5322_955_ngat) );
INVXL U_g3676 (.A(G4900_1093_gat), .Y(G4900_1093_ngat) );
INVXL U_g3677 (.A(G4903_671_gat), .Y(G4903_671_ngat) );
INVXL U_g3678 (.A(G5210_1094_gat), .Y(G5210_1094_ngat) );
INVXL U_g3679 (.A(G5213_672_gat), .Y(G5213_672_ngat) );
INVXL U_g3680 (.A(G7249_1024_gat), .Y(G7249_1024_ngat) );
INVXL U_g3681 (.A(G7256_1022_gat), .Y(G7256_1022_ngat) );
INVXL U_g3682 (.A(G3210_1026_gat), .Y(G3210_1026_ngat) );
INVXL U_g3683 (.A(G3211_827_gat), .Y(G3211_827_ngat) );
INVXL U_g3684 (.A(G5242_917_gat), .Y(G5242_917_ngat) );
INVXL U_g3685 (.A(G5245_830_gat), .Y(G5245_830_ngat) );
INVXL U_g3686 (.A(G5234_918_gat), .Y(G5234_918_ngat) );
INVXL U_g3687 (.A(G5237_720_gat), .Y(G5237_720_ngat) );
INVXL U_g3688 (.A(G5305_845_gat), .Y(G5305_845_ngat) );
INVXL U_g3689 (.A(G5312_1061_gat), .Y(G5312_1061_ngat) );
INVXL U_g3690 (.A(G5308_846_gat), .Y(G5308_846_ngat) );
INVXL U_g3691 (.A(G5311_1060_gat), .Y(G5311_1060_ngat) );
INVXL U_g3692 (.A(G5271_863_gat), .Y(G5271_863_ngat) );
INVXL U_g3693 (.A(G5278_1103_gat), .Y(G5278_1103_ngat) );
INVXL U_g3694 (.A(G5274_864_gat), .Y(G5274_864_ngat) );
INVXL U_g3695 (.A(G5277_1102_gat), .Y(G5277_1102_ngat) );
INVXL U_g3696 (.A(G6856_1327_gat), .Y(G6856_1327_ngat) );
INVXL U_g3697 (.A(G6859_431_gat), .Y(G6859_431_ngat) );
INVXL U_g3698 (.A(G6570_1329_gat), .Y(G6570_1329_ngat) );
INVXL U_g3699 (.A(G6573_432_gat), .Y(G6573_432_ngat) );
INVXL U_g3700 (.A(G6578_1350_gat), .Y(G6578_1350_ngat) );
INVXL U_g3701 (.A(G6581_433_gat), .Y(G6581_433_ngat) );
INVXL U_g3702 (.A(G6864_1352_gat), .Y(G6864_1352_ngat) );
INVXL U_g3703 (.A(G6867_434_gat), .Y(G6867_434_ngat) );
INVXL U_g3704 (.A(G6586_1378_gat), .Y(G6586_1378_ngat) );
INVXL U_g3705 (.A(G6589_435_gat), .Y(G6589_435_ngat) );
INVXL U_g3706 (.A(G6872_1377_gat), .Y(G6872_1377_ngat) );
INVXL U_g3707 (.A(G6875_436_gat), .Y(G6875_436_ngat) );
INVXL U_g3708 (.A(G6912_1374_gat), .Y(G6912_1374_ngat) );
INVXL U_g3709 (.A(G6915_437_gat), .Y(G6915_437_ngat) );
INVXL U_g3710 (.A(G6594_1375_gat), .Y(G6594_1375_ngat) );
INVXL U_g3711 (.A(G6597_438_gat), .Y(G6597_438_ngat) );
INVXL U_g3712 (.A(G6880_1361_gat), .Y(G6880_1361_ngat) );
INVXL U_g3713 (.A(G6883_439_gat), .Y(G6883_439_ngat) );
INVXL U_g3714 (.A(G6602_1359_gat), .Y(G6602_1359_ngat) );
INVXL U_g3715 (.A(G6605_440_gat), .Y(G6605_440_ngat) );
INVXL U_g3716 (.A(G6610_1266_gat), .Y(G6610_1266_ngat) );
INVXL U_g3717 (.A(G6613_441_gat), .Y(G6613_441_ngat) );
INVXL U_g3718 (.A(G6888_1267_gat), .Y(G6888_1267_ngat) );
INVXL U_g3719 (.A(G6891_442_gat), .Y(G6891_442_ngat) );
INVXL U_g3720 (.A(G6896_1302_gat), .Y(G6896_1302_ngat) );
INVXL U_g3721 (.A(G6899_443_gat), .Y(G6899_443_ngat) );
INVXL U_g3722 (.A(G6618_1303_gat), .Y(G6618_1303_ngat) );
INVXL U_g3723 (.A(G6621_444_gat), .Y(G6621_444_ngat) );
INVXL U_g3724 (.A(G6904_1296_gat), .Y(G6904_1296_ngat) );
INVXL U_g3725 (.A(G6907_445_gat), .Y(G6907_445_ngat) );
INVXL U_g3726 (.A(G6626_1297_gat), .Y(G6626_1297_ngat) );
INVXL U_g3727 (.A(G6629_446_gat), .Y(G6629_446_ngat) );
INVXL U_g3728 (.A(G6634_1275_gat), .Y(G6634_1275_ngat) );
INVXL U_g3729 (.A(G6637_447_gat), .Y(G6637_447_ngat) );
INVXL U_g3730 (.A(G6920_1276_gat), .Y(G6920_1276_ngat) );
INVXL U_g3731 (.A(G6923_448_gat), .Y(G6923_448_ngat) );
INVXL U_g3732 (.A(G5988_1290_gat), .Y(G5988_1290_ngat) );
INVXL U_g3733 (.A(G5991_449_gat), .Y(G5991_449_ngat) );
INVXL U_g3734 (.A(G5868_1291_gat), .Y(G5868_1291_ngat) );
INVXL U_g3735 (.A(G5871_450_gat), .Y(G5871_450_ngat) );
INVXL U_g3736 (.A(G5876_1259_gat), .Y(G5876_1259_ngat) );
INVXL U_g3737 (.A(G5879_451_gat), .Y(G5879_451_ngat) );
INVXL U_g3738 (.A(G5996_1260_gat), .Y(G5996_1260_ngat) );
INVXL U_g3739 (.A(G5999_452_gat), .Y(G5999_452_ngat) );
INVXL U_g3740 (.A(G6004_1254_gat), .Y(G6004_1254_ngat) );
INVXL U_g3741 (.A(G6007_453_gat), .Y(G6007_453_ngat) );
INVXL U_g3742 (.A(G5884_1255_gat), .Y(G5884_1255_ngat) );
INVXL U_g3743 (.A(G5887_454_gat), .Y(G5887_454_ngat) );
INVXL U_g3744 (.A(G6044_1251_gat), .Y(G6044_1251_ngat) );
INVXL U_g3745 (.A(G6047_455_gat), .Y(G6047_455_ngat) );
INVXL U_g3746 (.A(G5892_1250_gat), .Y(G5892_1250_ngat) );
INVXL U_g3747 (.A(G5895_456_gat), .Y(G5895_456_ngat) );
INVXL U_g3748 (.A(G5900_1288_gat), .Y(G5900_1288_ngat) );
INVXL U_g3749 (.A(G5903_457_gat), .Y(G5903_457_ngat) );
INVXL U_g3750 (.A(G6012_1287_gat), .Y(G6012_1287_ngat) );
INVXL U_g3751 (.A(G6015_458_gat), .Y(G6015_458_ngat) );
INVXL U_g3752 (.A(G6020_1395_gat), .Y(G6020_1395_ngat) );
INVXL U_g3753 (.A(G6023_459_gat), .Y(G6023_459_ngat) );
INVXL U_g3754 (.A(G5908_1394_gat), .Y(G5908_1394_ngat) );
INVXL U_g3755 (.A(G5911_460_gat), .Y(G5911_460_ngat) );
INVXL U_g3756 (.A(G5916_1390_gat), .Y(G5916_1390_ngat) );
INVXL U_g3757 (.A(G5919_461_gat), .Y(G5919_461_ngat) );
INVXL U_g3758 (.A(G6028_1389_gat), .Y(G6028_1389_ngat) );
INVXL U_g3759 (.A(G6031_462_gat), .Y(G6031_462_ngat) );
INVXL U_g3760 (.A(G6036_1383_gat), .Y(G6036_1383_ngat) );
INVXL U_g3761 (.A(G6039_463_gat), .Y(G6039_463_ngat) );
INVXL U_g3762 (.A(G5924_1382_gat), .Y(G5924_1382_ngat) );
INVXL U_g3763 (.A(G5927_464_gat), .Y(G5927_464_ngat) );
INVXL U_g3764 (.A(G7497_868_gat), .Y(G7497_868_ngat) );
INVXL U_g3765 (.A(G7504_1150_gat), .Y(G7504_1150_ngat) );
INVXL U_g3766 (.A(G6367_869_gat), .Y(G6367_869_ngat) );
INVXL U_g3767 (.A(G6374_1420_gat), .Y(G6374_1420_ngat) );
INVXL U_g3768 (.A(G5393_352_gat), .Y(G5393_352_ngat) );
INVXL U_g3769 (.A(G5400_1439_gat), .Y(G5400_1439_ngat) );
INVXL U_g3770 (.A(G5745_353_gat), .Y(G5745_353_ngat) );
INVXL U_g3771 (.A(G5752_1440_gat), .Y(G5752_1440_ngat) );
INVXL U_g3772 (.A(G7500_873_gat), .Y(G7500_873_ngat) );
INVXL U_g3773 (.A(G7503_1146_gat), .Y(G7503_1146_ngat) );
INVXL U_g3774 (.A(G6375_874_gat), .Y(G6375_874_ngat) );
INVXL U_g3775 (.A(G6382_1421_gat), .Y(G6382_1421_ngat) );
INVXL U_g3776 (.A(G5753_354_gat), .Y(G5753_354_ngat) );
INVXL U_g3777 (.A(G5760_1441_gat), .Y(G5760_1441_ngat) );
INVXL U_g3778 (.A(G5401_355_gat), .Y(G5401_355_ngat) );
INVXL U_g3779 (.A(G5408_1442_gat), .Y(G5408_1442_ngat) );
INVXL U_g3780 (.A(G6383_880_gat), .Y(G6383_880_ngat) );
INVXL U_g3781 (.A(G6390_1424_gat), .Y(G6390_1424_ngat) );
INVXL U_g3782 (.A(G7487_881_gat), .Y(G7487_881_ngat) );
INVXL U_g3783 (.A(G7494_1164_gat), .Y(G7494_1164_ngat) );
INVXL U_g3784 (.A(G5409_356_gat), .Y(G5409_356_ngat) );
INVXL U_g3785 (.A(G5416_1431_gat), .Y(G5416_1431_ngat) );
INVXL U_g3786 (.A(G5761_357_gat), .Y(G5761_357_ngat) );
INVXL U_g3787 (.A(G5768_1430_gat), .Y(G5768_1430_ngat) );
INVXL U_g3788 (.A(G5769_358_gat), .Y(G5769_358_ngat) );
INVXL U_g3789 (.A(G5776_1433_gat), .Y(G5776_1433_ngat) );
INVXL U_g3790 (.A(G5449_359_gat), .Y(G5449_359_ngat) );
INVXL U_g3791 (.A(G5456_1432_gat), .Y(G5456_1432_ngat) );
INVXL U_g3792 (.A(G7490_887_gat), .Y(G7490_887_ngat) );
INVXL U_g3793 (.A(G7493_1155_gat), .Y(G7493_1155_ngat) );
INVXL U_g3794 (.A(G6423_888_gat), .Y(G6423_888_ngat) );
INVXL U_g3795 (.A(G6430_1425_gat), .Y(G6430_1425_ngat) );
INVXL U_g3796 (.A(G7479_890_gat), .Y(G7479_890_ngat) );
INVXL U_g3797 (.A(G7486_1173_gat), .Y(G7486_1173_ngat) );
INVXL U_g3798 (.A(G6391_891_gat), .Y(G6391_891_ngat) );
INVXL U_g3799 (.A(G6398_1428_gat), .Y(G6398_1428_ngat) );
INVXL U_g3800 (.A(G5417_360_gat), .Y(G5417_360_ngat) );
INVXL U_g3801 (.A(G5424_1437_gat), .Y(G5424_1437_ngat) );
INVXL U_g3802 (.A(G5777_361_gat), .Y(G5777_361_ngat) );
INVXL U_g3803 (.A(G5784_1436_gat), .Y(G5784_1436_ngat) );
INVXL U_g3804 (.A(G5785_362_gat), .Y(G5785_362_ngat) );
INVXL U_g3805 (.A(G5792_1243_gat), .Y(G5792_1243_ngat) );
INVXL U_g3806 (.A(G5425_363_gat), .Y(G5425_363_ngat) );
INVXL U_g3807 (.A(G5432_1242_gat), .Y(G5432_1242_ngat) );
INVXL U_g3808 (.A(G6399_897_gat), .Y(G6399_897_ngat) );
INVXL U_g3809 (.A(G6406_1230_gat), .Y(G6406_1230_ngat) );
INVXL U_g3810 (.A(G7482_898_gat), .Y(G7482_898_ngat) );
INVXL U_g3811 (.A(G7485_1166_gat), .Y(G7485_1166_ngat) );
INVXL U_g3812 (.A(G7471_902_gat), .Y(G7471_902_ngat) );
INVXL U_g3813 (.A(G7478_1181_gat), .Y(G7478_1181_ngat) );
INVXL U_g3814 (.A(G6407_903_gat), .Y(G6407_903_ngat) );
INVXL U_g3815 (.A(G6414_1229_gat), .Y(G6414_1229_ngat) );
INVXL U_g3816 (.A(G5433_364_gat), .Y(G5433_364_ngat) );
INVXL U_g3817 (.A(G5440_1240_gat), .Y(G5440_1240_ngat) );
INVXL U_g3818 (.A(G5793_365_gat), .Y(G5793_365_ngat) );
INVXL U_g3819 (.A(G5800_1239_gat), .Y(G5800_1239_ngat) );
INVXL U_g3820 (.A(G5801_366_gat), .Y(G5801_366_ngat) );
INVXL U_g3821 (.A(G5808_1237_gat), .Y(G5808_1237_ngat) );
INVXL U_g3822 (.A(G5441_367_gat), .Y(G5441_367_ngat) );
INVXL U_g3823 (.A(G5448_1236_gat), .Y(G5448_1236_ngat) );
INVXL U_g3824 (.A(G6415_907_gat), .Y(G6415_907_ngat) );
INVXL U_g3825 (.A(G6422_1226_gat), .Y(G6422_1226_ngat) );
INVXL U_g3826 (.A(G7474_908_gat), .Y(G7474_908_ngat) );
INVXL U_g3827 (.A(G7477_1174_gat), .Y(G7477_1174_ngat) );
INVXL U_g3828 (.A(G5457_368_gat), .Y(G5457_368_ngat) );
INVXL U_g3829 (.A(G5464_1246_gat), .Y(G5464_1246_ngat) );
INVXL U_g3830 (.A(G6431_914_gat), .Y(G6431_914_ngat) );
INVXL U_g3831 (.A(G6438_1233_gat), .Y(G6438_1233_ngat) );
INVXL U_g3832 (.A(G5809_369_gat), .Y(G5809_369_ngat) );
INVXL U_g3833 (.A(G5816_1245_gat), .Y(G5816_1245_ngat) );
INVXL U_g3834 (.A(G7466_771_gat), .Y(G7466_771_ngat) );
INVXL U_g3835 (.A(G7469_1186_gat), .Y(G7469_1186_ngat) );
INVXL U_g3836 (.A(G6719_1202_gat), .Y(G6719_1202_ngat) );
INVXL U_g3837 (.A(G6720_1189_gat), .Y(G6720_1189_ngat) );
INVXL U_g3838 (.A(G6703_927_gat), .Y(G6703_927_ngat) );
INVXL U_g3839 (.A(G6710_1213_gat), .Y(G6710_1213_ngat) );
INVXL U_g3840 (.A(G6519_928_gat), .Y(G6519_928_ngat) );
INVXL U_g3841 (.A(G6526_1418_gat), .Y(G6526_1418_ngat) );
INVXL U_g3842 (.A(G4881_375_gat), .Y(G4881_375_ngat) );
INVXL U_g3843 (.A(G4888_1460_gat), .Y(G4888_1460_ngat) );
INVXL U_g3844 (.A(G5191_376_gat), .Y(G5191_376_ngat) );
INVXL U_g3845 (.A(G5198_1461_gat), .Y(G5198_1461_ngat) );
INVXL U_g3846 (.A(G5199_377_gat), .Y(G5199_377_ngat) );
INVXL U_g3847 (.A(G5206_1444_gat), .Y(G5206_1444_ngat) );
INVXL U_g3848 (.A(G4889_378_gat), .Y(G4889_378_ngat) );
INVXL U_g3849 (.A(G4896_1445_gat), .Y(G4896_1445_ngat) );
INVXL U_g3850 (.A(G6527_932_gat), .Y(G6527_932_ngat) );
INVXL U_g3851 (.A(G6534_1408_gat), .Y(G6534_1408_ngat) );
INVXL U_g3852 (.A(G6706_933_gat), .Y(G6706_933_ngat) );
INVXL U_g3853 (.A(G6709_1206_gat), .Y(G6709_1206_ngat) );
INVXL U_g3854 (.A(G5215_379_gat), .Y(G5215_379_ngat) );
INVXL U_g3855 (.A(G5222_1450_gat), .Y(G5222_1450_ngat) );
INVXL U_g3856 (.A(G6543_937_gat), .Y(G6543_937_ngat) );
INVXL U_g3857 (.A(G6550_1412_gat), .Y(G6550_1412_ngat) );
INVXL U_g3858 (.A(G6698_938_gat), .Y(G6698_938_ngat) );
INVXL U_g3859 (.A(G6701_1281_gat), .Y(G6701_1281_ngat) );
INVXL U_g3860 (.A(G4905_380_gat), .Y(G4905_380_ngat) );
INVXL U_g3861 (.A(G4912_1451_gat), .Y(G4912_1451_ngat) );
INVXL U_g3862 (.A(G4921_381_gat), .Y(G4921_381_ngat) );
INVXL U_g3863 (.A(G4928_1454_gat), .Y(G4928_1454_ngat) );
INVXL U_g3864 (.A(G6559_944_gat), .Y(G6559_944_ngat) );
INVXL U_g3865 (.A(G6566_1414_gat), .Y(G6566_1414_ngat) );
INVXL U_g3866 (.A(G5223_382_gat), .Y(G5223_382_ngat) );
INVXL U_g3867 (.A(G5230_1455_gat), .Y(G5230_1455_ngat) );
INVXL U_g3868 (.A(G6690_780_gat), .Y(G6690_780_ngat) );
INVXL U_g3869 (.A(G6693_1222_gat), .Y(G6693_1222_ngat) );
INVXL U_g3870 (.A(G7296_811_gat), .Y(G7296_811_ngat) );
INVXL U_g3871 (.A(G7299_1232_gat), .Y(G7299_1232_ngat) );
INVXL U_g3872 (.A(G6418_947_gat), .Y(G6418_947_ngat) );
INVXL U_g3873 (.A(G6421_1180_gat), .Y(G6421_1180_ngat) );
INVXL U_g3874 (.A(G7304_948_gat), .Y(G7304_948_ngat) );
INVXL U_g3875 (.A(G7307_1228_gat), .Y(G7307_1228_ngat) );
INVXL U_g3876 (.A(G7301_949_gat), .Y(G7301_949_ngat) );
INVXL U_g3877 (.A(G7308_1227_gat), .Y(G7308_1227_ngat) );
INVXL U_g3878 (.A(G6410_950_gat), .Y(G6410_950_ngat) );
INVXL U_g3879 (.A(G6413_1175_gat), .Y(G6413_1175_ngat) );
INVXL U_g3880 (.A(G6402_951_gat), .Y(G6402_951_ngat) );
INVXL U_g3881 (.A(G6405_1172_gat), .Y(G6405_1172_ngat) );
INVXL U_g3882 (.A(G7312_952_gat), .Y(G7312_952_ngat) );
INVXL U_g3883 (.A(G7315_1427_gat), .Y(G7315_1427_ngat) );
INVXL U_g3884 (.A(G6434_954_gat), .Y(G6434_954_ngat) );
INVXL U_g3885 (.A(G6437_1187_gat), .Y(G6437_1187_ngat) );
INVXL U_g3886 (.A(G5318_816_gat), .Y(G5318_816_ngat) );
INVXL U_g3887 (.A(G5321_1244_gat), .Y(G5321_1244_ngat) );
INVXL U_g3888 (.A(G5326_956_gat), .Y(G5326_956_ngat) );
INVXL U_g3889 (.A(G5329_1238_gat), .Y(G5329_1238_ngat) );
INVXL U_g3890 (.A(G5323_959_gat), .Y(G5323_959_ngat) );
INVXL U_g3891 (.A(G5330_1235_gat), .Y(G5330_1235_ngat) );
INVXL U_g3892 (.A(G5334_962_gat), .Y(G5334_962_ngat) );
INVXL U_g3893 (.A(G5337_1435_gat), .Y(G5337_1435_ngat) );
INVXL U_g3894 (.A(G7224_1270_gat), .Y(G7224_1270_ngat) );
INVXL U_g3895 (.A(G7227_1358_gat), .Y(G7227_1358_ngat) );
INVXL U_g3896 (.A(G7205_1273_gat), .Y(G7205_1273_ngat) );
INVXL U_g3897 (.A(G7212_1277_gat), .Y(G7212_1277_ngat) );
INVXL U_g3898 (.A(G6721_1274_gat), .Y(G6721_1274_ngat) );
INVXL U_g3899 (.A(G6728_1278_gat), .Y(G6728_1278_ngat) );
INVXL U_g3900 (.A(G4897_548_gat), .Y(G4897_548_ngat) );
INVXL U_g3901 (.A(G4904_1448_gat), .Y(G4904_1448_ngat) );
INVXL U_g3902 (.A(G5207_549_gat), .Y(G5207_549_ngat) );
INVXL U_g3903 (.A(G5214_1449_gat), .Y(G5214_1449_ngat) );
INVXL U_g3904 (.A(G6695_983_gat), .Y(G6695_983_ngat) );
INVXL U_g3905 (.A(G6702_1216_gat), .Y(G6702_1216_ngat) );
INVXL U_g3906 (.A(G6535_984_gat), .Y(G6535_984_ngat) );
INVXL U_g3907 (.A(G6542_1410_gat), .Y(G6542_1410_ngat) );
INVXL U_g3908 (.A(G7265_1285_gat), .Y(G7265_1285_ngat) );
INVXL U_g3909 (.A(G7272_1399_gat), .Y(G7272_1399_ngat) );
INVXL U_g3910 (.A(G6463_1309_gat), .Y(G6463_1309_ngat) );
INVXL U_g3911 (.A(G6470_1357_gat), .Y(G6470_1357_ngat) );
INVXL U_g3912 (.A(G6495_1311_gat), .Y(G6495_1311_ngat) );
INVXL U_g3913 (.A(G6502_1371_gat), .Y(G6502_1371_ngat) );
INVXL U_g3914 (.A(G7551_1316_gat), .Y(G7551_1316_ngat) );
INVXL U_g3915 (.A(G7558_1341_gat), .Y(G7558_1341_ngat) );
INVXL U_g3916 (.A(G7401_1318_gat), .Y(G7401_1318_ngat) );
INVXL U_g3917 (.A(G7408_1391_gat), .Y(G7408_1391_ngat) );
INVXL U_g3918 (.A(G7393_1319_gat), .Y(G7393_1319_ngat) );
INVXL U_g3919 (.A(G7400_1398_gat), .Y(G7400_1398_ngat) );
INVXL U_g3920 (.A(G7409_1321_gat), .Y(G7409_1321_ngat) );
INVXL U_g3921 (.A(G7416_1386_gat), .Y(G7416_1386_ngat) );
INVXL U_g3922 (.A(G7507_1002_gat), .Y(G7507_1002_ngat) );
INVXL U_g3923 (.A(G7514_1326_gat), .Y(G7514_1326_ngat) );
INVXL U_g3924 (.A(G7510_1003_gat), .Y(G7510_1003_ngat) );
INVXL U_g3925 (.A(G7513_1325_gat), .Y(G7513_1325_ngat) );
INVXL U_g3926 (.A(G7239_1005_gat), .Y(G7239_1005_ngat) );
INVXL U_g3927 (.A(G7246_1355_gat), .Y(G7246_1355_ngat) );
INVXL U_g3928 (.A(G6439_1333_gat), .Y(G6439_1333_ngat) );
INVXL U_g3929 (.A(G6446_1332_gat), .Y(G6446_1332_ngat) );
INVXL U_g3930 (.A(G6447_1335_gat), .Y(G6447_1335_ngat) );
INVXL U_g3931 (.A(G6454_1354_gat), .Y(G6454_1354_ngat) );
INVXL U_g3932 (.A(G6455_1337_gat), .Y(G6455_1337_ngat) );
INVXL U_g3933 (.A(G6462_1380_gat), .Y(G6462_1380_ngat) );
INVXL U_g3934 (.A(G7242_1018_gat), .Y(G7242_1018_ngat) );
INVXL U_g3935 (.A(G7245_1331_gat), .Y(G7245_1331_ngat) );
INVXL U_g3936 (.A(G7252_825_gat), .Y(G7252_825_ngat) );
INVXL U_g3937 (.A(G7255_1364_gat), .Y(G7255_1364_ngat) );
INVXL U_g3938 (.A(G6765_1365_gat), .Y(G6765_1365_ngat) );
INVXL U_g3939 (.A(G6772_1363_gat), .Y(G6772_1363_ngat) );
INVXL U_g3940 (.A(G5239_719_gat), .Y(G5239_719_ngat) );
INVXL U_g3941 (.A(G5246_1194_gat), .Y(G5246_1194_ngat) );
INVXL U_g3942 (.A(G5231_561_gat), .Y(G5231_561_ngat) );
INVXL U_g3943 (.A(G5238_1195_gat), .Y(G5238_1195_ngat) );
INVXL U_g3944 (.A(G7232_1033_gat), .Y(G7232_1033_ngat) );
INVXL U_g3945 (.A(G7235_1381_gat), .Y(G7235_1381_ngat) );
INVXL U_g3946 (.A(G7229_1037_gat), .Y(G7229_1037_ngat) );
INVXL U_g3947 (.A(G7236_1372_gat), .Y(G7236_1372_ngat) );
INVXL U_g3948 (.A(G7260_1040_gat), .Y(G7260_1040_ngat) );
INVXL U_g3949 (.A(G7263_1393_gat), .Y(G7263_1393_ngat) );
INVXL U_g3950 (.A(G7257_1043_gat), .Y(G7257_1043_ngat) );
INVXL U_g3951 (.A(G7264_1387_gat), .Y(G7264_1387_ngat) );
INVXL U_g3952 (.A(G7428_1404_gat), .Y(G7428_1404_ngat) );
INVXL U_g3953 (.A(G7431_1401_gat), .Y(G7431_1401_ngat) );
INVXL U_g3954 (.A(G3682_839_gat), .Y(G3682_839_ngat) );
INVXL U_g3955 (.A(G4389_1405_gat), .Y(G4389_1405_ngat) );
INVXL U_g3956 (.A(G5284_1051_gat), .Y(G5284_1051_ngat) );
INVXL U_g3957 (.A(G5287_1413_gat), .Y(G5287_1413_ngat) );
INVXL U_g3958 (.A(G5300_1052_gat), .Y(G5300_1052_ngat) );
INVXL U_g3959 (.A(G5303_1417_gat), .Y(G5303_1417_ngat) );
INVXL U_g3960 (.A(G6530_1053_gat), .Y(G6530_1053_ngat) );
INVXL U_g3961 (.A(G6533_1212_gat), .Y(G6533_1212_ngat) );
INVXL U_g3962 (.A(G5289_1054_gat), .Y(G5289_1054_ngat) );
INVXL U_g3963 (.A(G5296_1411_gat), .Y(G5296_1411_ngat) );
INVXL U_g3964 (.A(G6538_1055_gat), .Y(G6538_1055_ngat) );
INVXL U_g3965 (.A(G6541_1282_gat), .Y(G6541_1282_ngat) );
INVXL U_g3966 (.A(G5292_1056_gat), .Y(G5292_1056_ngat) );
INVXL U_g3967 (.A(G5295_1409_gat), .Y(G5295_1409_ngat) );
INVXL U_g3968 (.A(G6546_1057_gat), .Y(G6546_1057_ngat) );
INVXL U_g3969 (.A(G6549_1215_gat), .Y(G6549_1215_ngat) );
INVXL U_g3970 (.A(G5281_1058_gat), .Y(G5281_1058_ngat) );
INVXL U_g3971 (.A(G5288_1406_gat), .Y(G5288_1406_ngat) );
INVXL U_g3972 (.A(G6562_1059_gat), .Y(G6562_1059_ngat) );
INVXL U_g3973 (.A(G6565_1223_gat), .Y(G6565_1223_ngat) );
INVXL U_g3974 (.A(G5313_1416_gat), .Y(G5313_1416_ngat) );
INVXL U_g3975 (.A(G5314_1415_gat), .Y(G5314_1415_ngat) );
INVXL U_g3976 (.A(G5297_1062_gat), .Y(G5297_1062_ngat) );
INVXL U_g3977 (.A(G5304_1407_gat), .Y(G5304_1407_ngat) );
INVXL U_g3978 (.A(G6522_1063_gat), .Y(G6522_1063_ngat) );
INVXL U_g3979 (.A(G6525_1207_gat), .Y(G6525_1207_ngat) );
INVXL U_g3980 (.A(G7327_1064_gat), .Y(G7327_1064_ngat) );
INVXL U_g3981 (.A(G7334_1422_gat), .Y(G7334_1422_ngat) );
INVXL U_g3982 (.A(G6370_1065_gat), .Y(G6370_1065_ngat) );
INVXL U_g3983 (.A(G6373_1147_gat), .Y(G6373_1147_ngat) );
INVXL U_g3984 (.A(G6378_1066_gat), .Y(G6378_1066_ngat) );
INVXL U_g3985 (.A(G6381_1151_gat), .Y(G6381_1151_ngat) );
INVXL U_g3986 (.A(G7330_1067_gat), .Y(G7330_1067_ngat) );
INVXL U_g3987 (.A(G7333_1419_gat), .Y(G7333_1419_ngat) );
INVXL U_g3988 (.A(G7317_1068_gat), .Y(G7317_1068_ngat) );
INVXL U_g3989 (.A(G7324_1426_gat), .Y(G7324_1426_ngat) );
INVXL U_g3990 (.A(G6386_1069_gat), .Y(G6386_1069_ngat) );
INVXL U_g3991 (.A(G6389_1154_gat), .Y(G6389_1154_ngat) );
INVXL U_g3992 (.A(G6426_1070_gat), .Y(G6426_1070_ngat) );
INVXL U_g3993 (.A(G6429_1165_gat), .Y(G6429_1165_ngat) );
INVXL U_g3994 (.A(G7320_1071_gat), .Y(G7320_1071_ngat) );
INVXL U_g3995 (.A(G7323_1423_gat), .Y(G7323_1423_ngat) );
INVXL U_g3996 (.A(G7309_1072_gat), .Y(G7309_1072_ngat) );
INVXL U_g3997 (.A(G7316_1231_gat), .Y(G7316_1231_ngat) );
INVXL U_g3998 (.A(G6394_1073_gat), .Y(G6394_1073_ngat) );
INVXL U_g3999 (.A(G6397_1167_gat), .Y(G6397_1167_ngat) );
INVXL U_g4000 (.A(G5339_1074_gat), .Y(G5339_1074_ngat) );
INVXL U_g4001 (.A(G5346_1434_gat), .Y(G5346_1434_ngat) );
INVXL U_g4002 (.A(G5342_1079_gat), .Y(G5342_1079_ngat) );
INVXL U_g4003 (.A(G5345_1429_gat), .Y(G5345_1429_ngat) );
INVXL U_g4004 (.A(G5331_1080_gat), .Y(G5331_1080_ngat) );
INVXL U_g4005 (.A(G5338_1241_gat), .Y(G5338_1241_ngat) );
INVXL U_g4006 (.A(G5349_1083_gat), .Y(G5349_1083_ngat) );
INVXL U_g4007 (.A(G5356_1443_gat), .Y(G5356_1443_ngat) );
INVXL U_g4008 (.A(G5352_1088_gat), .Y(G5352_1088_ngat) );
INVXL U_g4009 (.A(G5355_1438_gat), .Y(G5355_1438_ngat) );
INVXL U_g4010 (.A(G5266_1091_gat), .Y(G5266_1091_ngat) );
INVXL U_g4011 (.A(G5269_1459_gat), .Y(G5269_1459_ngat) );
INVXL U_g4012 (.A(G5255_1092_gat), .Y(G5255_1092_ngat) );
INVXL U_g4013 (.A(G5262_1452_gat), .Y(G5262_1452_ngat) );
INVXL U_g4014 (.A(G5258_1097_gat), .Y(G5258_1097_ngat) );
INVXL U_g4015 (.A(G5261_1447_gat), .Y(G5261_1447_ngat) );
INVXL U_g4016 (.A(G5247_1098_gat), .Y(G5247_1098_ngat) );
INVXL U_g4017 (.A(G5254_1456_gat), .Y(G5254_1456_ngat) );
INVXL U_g4018 (.A(G5250_1101_gat), .Y(G5250_1101_ngat) );
INVXL U_g4019 (.A(G5253_1453_gat), .Y(G5253_1453_ngat) );
INVXL U_g4020 (.A(G5279_1458_gat), .Y(G5279_1458_ngat) );
INVXL U_g4021 (.A(G5280_1457_gat), .Y(G5280_1457_ngat) );
INVXL U_g4022 (.A(G5263_1104_gat), .Y(G5263_1104_ngat) );
INVXL U_g4023 (.A(G5270_1446_gat), .Y(G5270_1446_ngat) );
INVXL U_g4024 (.A(G6853_318_gat), .Y(G6853_318_ngat) );
INVXL U_g4025 (.A(G6860_1665_gat), .Y(G6860_1665_ngat) );
INVXL U_g4026 (.A(G6567_319_gat), .Y(G6567_319_ngat) );
INVXL U_g4027 (.A(G6574_1667_gat), .Y(G6574_1667_ngat) );
INVXL U_g4028 (.A(G6575_320_gat), .Y(G6575_320_ngat) );
INVXL U_g4029 (.A(G6582_1688_gat), .Y(G6582_1688_ngat) );
INVXL U_g4030 (.A(G6861_321_gat), .Y(G6861_321_ngat) );
INVXL U_g4031 (.A(G6868_1690_gat), .Y(G6868_1690_ngat) );
INVXL U_g4032 (.A(G6583_322_gat), .Y(G6583_322_ngat) );
INVXL U_g4033 (.A(G6590_1707_gat), .Y(G6590_1707_ngat) );
INVXL U_g4034 (.A(G6869_323_gat), .Y(G6869_323_ngat) );
INVXL U_g4035 (.A(G6876_1706_gat), .Y(G6876_1706_ngat) );
INVXL U_g4036 (.A(G6909_324_gat), .Y(G6909_324_ngat) );
INVXL U_g4037 (.A(G6916_1703_gat), .Y(G6916_1703_ngat) );
INVXL U_g4038 (.A(G6591_325_gat), .Y(G6591_325_ngat) );
INVXL U_g4039 (.A(G6598_1704_gat), .Y(G6598_1704_ngat) );
INVXL U_g4040 (.A(G6877_326_gat), .Y(G6877_326_ngat) );
INVXL U_g4041 (.A(G6884_1694_gat), .Y(G6884_1694_ngat) );
INVXL U_g4042 (.A(G6599_327_gat), .Y(G6599_327_ngat) );
INVXL U_g4043 (.A(G6606_1692_gat), .Y(G6606_1692_ngat) );
INVXL U_g4044 (.A(G6607_328_gat), .Y(G6607_328_ngat) );
INVXL U_g4045 (.A(G6614_1602_gat), .Y(G6614_1602_ngat) );
INVXL U_g4046 (.A(G6885_329_gat), .Y(G6885_329_ngat) );
INVXL U_g4047 (.A(G6892_1603_gat), .Y(G6892_1603_ngat) );
INVXL U_g4048 (.A(G6893_330_gat), .Y(G6893_330_ngat) );
INVXL U_g4049 (.A(G6900_1635_gat), .Y(G6900_1635_ngat) );
INVXL U_g4050 (.A(G6615_331_gat), .Y(G6615_331_ngat) );
INVXL U_g4051 (.A(G6622_1636_gat), .Y(G6622_1636_ngat) );
INVXL U_g4052 (.A(G6901_332_gat), .Y(G6901_332_ngat) );
INVXL U_g4053 (.A(G6908_1630_gat), .Y(G6908_1630_ngat) );
INVXL U_g4054 (.A(G6623_333_gat), .Y(G6623_333_ngat) );
INVXL U_g4055 (.A(G6630_1631_gat), .Y(G6630_1631_ngat) );
INVXL U_g4056 (.A(G6631_334_gat), .Y(G6631_334_ngat) );
INVXL U_g4057 (.A(G6638_1612_gat), .Y(G6638_1612_ngat) );
INVXL U_g4058 (.A(G6917_335_gat), .Y(G6917_335_ngat) );
INVXL U_g4059 (.A(G6924_1613_gat), .Y(G6924_1613_ngat) );
INVXL U_g4060 (.A(G5985_336_gat), .Y(G5985_336_ngat) );
INVXL U_g4061 (.A(G5992_1625_gat), .Y(G5992_1625_ngat) );
INVXL U_g4062 (.A(G5865_337_gat), .Y(G5865_337_ngat) );
INVXL U_g4063 (.A(G5872_1626_gat), .Y(G5872_1626_ngat) );
INVXL U_g4064 (.A(G5873_338_gat), .Y(G5873_338_ngat) );
INVXL U_g4065 (.A(G5880_1596_gat), .Y(G5880_1596_ngat) );
INVXL U_g4066 (.A(G5993_339_gat), .Y(G5993_339_ngat) );
INVXL U_g4067 (.A(G6000_1597_gat), .Y(G6000_1597_ngat) );
INVXL U_g4068 (.A(G6001_340_gat), .Y(G6001_340_ngat) );
INVXL U_g4069 (.A(G6008_1592_gat), .Y(G6008_1592_ngat) );
INVXL U_g4070 (.A(G5881_341_gat), .Y(G5881_341_ngat) );
INVXL U_g4071 (.A(G5888_1593_gat), .Y(G5888_1593_ngat) );
INVXL U_g4072 (.A(G6041_342_gat), .Y(G6041_342_ngat) );
INVXL U_g4073 (.A(G6048_1589_gat), .Y(G6048_1589_ngat) );
INVXL U_g4074 (.A(G5889_343_gat), .Y(G5889_343_ngat) );
INVXL U_g4075 (.A(G5896_1588_gat), .Y(G5896_1588_ngat) );
INVXL U_g4076 (.A(G5897_344_gat), .Y(G5897_344_ngat) );
INVXL U_g4077 (.A(G5904_1623_gat), .Y(G5904_1623_ngat) );
INVXL U_g4078 (.A(G6009_345_gat), .Y(G6009_345_ngat) );
INVXL U_g4079 (.A(G6016_1622_gat), .Y(G6016_1622_ngat) );
INVXL U_g4080 (.A(G6017_346_gat), .Y(G6017_346_ngat) );
INVXL U_g4081 (.A(G6024_1718_gat), .Y(G6024_1718_ngat) );
INVXL U_g4082 (.A(G5905_347_gat), .Y(G5905_347_ngat) );
INVXL U_g4083 (.A(G5912_1717_gat), .Y(G5912_1717_ngat) );
INVXL U_g4084 (.A(G5913_348_gat), .Y(G5913_348_ngat) );
INVXL U_g4085 (.A(G5920_1715_gat), .Y(G5920_1715_ngat) );
INVXL U_g4086 (.A(G6025_349_gat), .Y(G6025_349_ngat) );
INVXL U_g4087 (.A(G6032_1714_gat), .Y(G6032_1714_ngat) );
INVXL U_g4088 (.A(G6033_350_gat), .Y(G6033_350_ngat) );
INVXL U_g4089 (.A(G6040_1710_gat), .Y(G6040_1710_ngat) );
INVXL U_g4090 (.A(G5921_351_gat), .Y(G5921_351_ngat) );
INVXL U_g4091 (.A(G5928_1709_gat), .Y(G5928_1709_ngat) );
INVXL U_g4092 (.A(G7505_1511_gat), .Y(G7505_1511_ngat) );
INVXL U_g4093 (.A(G7506_1507_gat), .Y(G7506_1507_ngat) );
INVXL U_g4094 (.A(G2954_1740_gat), .Y(G2954_1740_ngat) );
INVXL U_g4095 (.A(G2955_1508_gat), .Y(G2955_1508_ngat) );
INVXL U_g4096 (.A(G1544_1148_gat), .Y(G1544_1148_ngat) );
INVXL U_g4097 (.A(G1545_1509_gat), .Y(G1545_1509_ngat) );
INVXL U_g4098 (.A(G1793_1149_gat), .Y(G1793_1149_ngat) );
INVXL U_g4099 (.A(G1794_1510_gat), .Y(G1794_1510_ngat) );
INVXL U_g4100 (.A(G2963_1741_gat), .Y(G2963_1741_ngat) );
INVXL U_g4101 (.A(G2964_1512_gat), .Y(G2964_1512_ngat) );
INVXL U_g4102 (.A(G1803_1152_gat), .Y(G1803_1152_ngat) );
INVXL U_g4103 (.A(G1804_1513_gat), .Y(G1804_1513_ngat) );
INVXL U_g4104 (.A(G1554_1153_gat), .Y(G1554_1153_ngat) );
INVXL U_g4105 (.A(G1555_1514_gat), .Y(G1555_1514_ngat) );
INVXL U_g4106 (.A(G2971_1744_gat), .Y(G2971_1744_ngat) );
INVXL U_g4107 (.A(G2972_1515_gat), .Y(G2972_1515_ngat) );
INVXL U_g4108 (.A(G7495_1523_gat), .Y(G7495_1523_ngat) );
INVXL U_g4109 (.A(G7496_1516_gat), .Y(G7496_1516_ngat) );
INVXL U_g4110 (.A(G1571_1156_gat), .Y(G1571_1156_ngat) );
INVXL U_g4111 (.A(G1572_1517_gat), .Y(G1572_1517_ngat) );
INVXL U_g4112 (.A(G1820_1157_gat), .Y(G1820_1157_ngat) );
INVXL U_g4113 (.A(G1821_1518_gat), .Y(G1821_1518_ngat) );
INVXL U_g4114 (.A(G1848_1160_gat), .Y(G1848_1160_ngat) );
INVXL U_g4115 (.A(G1849_1521_gat), .Y(G1849_1521_ngat) );
INVXL U_g4116 (.A(G1685_1163_gat), .Y(G1685_1163_ngat) );
INVXL U_g4117 (.A(G1686_1522_gat), .Y(G1686_1522_ngat) );
INVXL U_g4118 (.A(G3016_1745_gat), .Y(G3016_1745_ngat) );
INVXL U_g4119 (.A(G3017_1524_gat), .Y(G3017_1524_ngat) );
INVXL U_g4120 (.A(G4547_1532_gat), .Y(G4547_1532_ngat) );
INVXL U_g4121 (.A(G4548_1525_gat), .Y(G4548_1525_ngat) );
INVXL U_g4122 (.A(G2980_1748_gat), .Y(G2980_1748_ngat) );
INVXL U_g4123 (.A(G2981_1526_gat), .Y(G2981_1526_ngat) );
INVXL U_g4124 (.A(G1596_1168_gat), .Y(G1596_1168_ngat) );
INVXL U_g4125 (.A(G1597_1527_gat), .Y(G1597_1527_ngat) );
INVXL U_g4126 (.A(G1857_1169_gat), .Y(G1857_1169_ngat) );
INVXL U_g4127 (.A(G1858_1528_gat), .Y(G1858_1528_ngat) );
INVXL U_g4128 (.A(G1867_1170_gat), .Y(G1867_1170_ngat) );
INVXL U_g4129 (.A(G1868_1529_gat), .Y(G1868_1529_ngat) );
INVXL U_g4130 (.A(G1607_1171_gat), .Y(G1607_1171_ngat) );
INVXL U_g4131 (.A(G1608_1530_gat), .Y(G1608_1530_ngat) );
INVXL U_g4132 (.A(G2990_1579_gat), .Y(G2990_1579_ngat) );
INVXL U_g4133 (.A(G2991_1531_gat), .Y(G2991_1531_ngat) );
INVXL U_g4134 (.A(G4538_1540_gat), .Y(G4538_1540_ngat) );
INVXL U_g4135 (.A(G4539_1533_gat), .Y(G4539_1533_ngat) );
INVXL U_g4136 (.A(G2999_1578_gat), .Y(G2999_1578_ngat) );
INVXL U_g4137 (.A(G3000_1534_gat), .Y(G3000_1534_ngat) );
INVXL U_g4138 (.A(G1628_1176_gat), .Y(G1628_1176_ngat) );
INVXL U_g4139 (.A(G1629_1535_gat), .Y(G1629_1535_ngat) );
INVXL U_g4140 (.A(G1883_1177_gat), .Y(G1883_1177_ngat) );
INVXL U_g4141 (.A(G1884_1536_gat), .Y(G1884_1536_ngat) );
INVXL U_g4142 (.A(G1901_1178_gat), .Y(G1901_1178_ngat) );
INVXL U_g4143 (.A(G1902_1537_gat), .Y(G1902_1537_ngat) );
INVXL U_g4144 (.A(G1653_1179_gat), .Y(G1653_1179_ngat) );
INVXL U_g4145 (.A(G1654_1538_gat), .Y(G1654_1538_ngat) );
INVXL U_g4146 (.A(G3007_1575_gat), .Y(G3007_1575_ngat) );
INVXL U_g4147 (.A(G3008_1539_gat), .Y(G3008_1539_ngat) );
INVXL U_g4148 (.A(G1693_1184_gat), .Y(G1693_1184_ngat) );
INVXL U_g4149 (.A(G1694_1542_gat), .Y(G1694_1542_ngat) );
INVXL U_g4150 (.A(G4529_1545_gat), .Y(G4529_1545_ngat) );
INVXL U_g4151 (.A(G4530_1185_gat), .Y(G4530_1185_ngat) );
INVXL U_g4152 (.A(G3019_1581_gat), .Y(G3019_1581_ngat) );
INVXL U_g4153 (.A(G3020_1543_gat), .Y(G3020_1543_ngat) );
INVXL U_g4154 (.A(G1919_1188_gat), .Y(G1919_1188_ngat) );
INVXL U_g4155 (.A(G1920_1544_gat), .Y(G1920_1544_ngat) );
INVXL U_g4156 (.A(G912_1550_gat), .Y(G912_1550_ngat) );
INVXL U_g4157 (.A(G906_1554_gat), .Y(G906_1554_ngat) );
INVXL U_g4158 (.A(G1121_1552_gat), .Y(G1121_1552_ngat) );
INVXL U_g4159 (.A(G1112_1553_gat), .Y(G1112_1553_ngat) );
INVXL U_g4160 (.A(G3520_1564_gat), .Y(G3520_1564_ngat) );
INVXL U_g4161 (.A(G3521_1557_gat), .Y(G3521_1557_ngat) );
INVXL U_g4162 (.A(G3174_1738_gat), .Y(G3174_1738_ngat) );
INVXL U_g4163 (.A(G3175_1558_gat), .Y(G3175_1558_ngat) );
INVXL U_g4164 (.A(G790_1208_gat), .Y(G790_1208_ngat) );
INVXL U_g4165 (.A(G791_1559_gat), .Y(G791_1559_ngat) );
INVXL U_g4166 (.A(G1024_1209_gat), .Y(G1024_1209_ngat) );
INVXL U_g4167 (.A(G1025_1560_gat), .Y(G1025_1560_ngat) );
INVXL U_g4168 (.A(G1036_1210_gat), .Y(G1036_1210_ngat) );
INVXL U_g4169 (.A(G1037_1561_gat), .Y(G1037_1561_ngat) );
INVXL U_g4170 (.A(G803_1211_gat), .Y(G803_1211_ngat) );
INVXL U_g4171 (.A(G804_1562_gat), .Y(G804_1562_ngat) );
INVXL U_g4172 (.A(G3184_1729_gat), .Y(G3184_1729_ngat) );
INVXL U_g4173 (.A(G3185_1563_gat), .Y(G3185_1563_ngat) );
INVXL U_g4174 (.A(G1072_1214_gat), .Y(G1072_1214_ngat) );
INVXL U_g4175 (.A(G1073_1565_gat), .Y(G1073_1565_ngat) );
INVXL U_g4176 (.A(G3201_1733_gat), .Y(G3201_1733_ngat) );
INVXL U_g4177 (.A(G3202_1566_gat), .Y(G3202_1566_ngat) );
INVXL U_g4178 (.A(G3511_1567_gat), .Y(G3511_1567_ngat) );
INVXL U_g4179 (.A(G3512_1616_gat), .Y(G3512_1616_ngat) );
INVXL U_g4180 (.A(G851_1217_gat), .Y(G851_1217_ngat) );
INVXL U_g4181 (.A(G852_1568_gat), .Y(G852_1568_ngat) );
INVXL U_g4182 (.A(G893_1220_gat), .Y(G893_1220_ngat) );
INVXL U_g4183 (.A(G894_1570_gat), .Y(G894_1570_ngat) );
INVXL U_g4184 (.A(G3502_1573_gat), .Y(G3502_1573_ngat) );
INVXL U_g4185 (.A(G3503_1221_gat), .Y(G3503_1221_ngat) );
INVXL U_g4186 (.A(G3213_1735_gat), .Y(G3213_1735_ngat) );
INVXL U_g4187 (.A(G3214_1571_gat), .Y(G3214_1571_ngat) );
INVXL U_g4188 (.A(G1091_1224_gat), .Y(G1091_1224_ngat) );
INVXL U_g4189 (.A(G1092_1572_gat), .Y(G1092_1572_ngat) );
INVXL U_g4190 (.A(G4224_1574_gat), .Y(G4224_1574_ngat) );
INVXL U_g4191 (.A(G4225_1225_gat), .Y(G4225_1225_ngat) );
INVXL U_g4192 (.A(G4233_1576_gat), .Y(G4233_1576_ngat) );
INVXL U_g4193 (.A(G4234_1577_gat), .Y(G4234_1577_ngat) );
INVXL U_g4194 (.A(G4242_1580_gat), .Y(G4242_1580_ngat) );
INVXL U_g4195 (.A(G4243_1747_gat), .Y(G4243_1747_ngat) );
INVXL U_g4196 (.A(G1261_1582_gat), .Y(G1261_1582_ngat) );
INVXL U_g4197 (.A(G1262_1234_gat), .Y(G1262_1234_ngat) );
INVXL U_g4198 (.A(G1270_1583_gat), .Y(G1270_1583_ngat) );
INVXL U_g4199 (.A(G1271_1584_gat), .Y(G1271_1584_ngat) );
INVXL U_g4200 (.A(G1279_1585_gat), .Y(G1279_1585_ngat) );
INVXL U_g4201 (.A(G1280_1751_gat), .Y(G1280_1751_ngat) );
INVXL U_g4202 (.A(G7276_1247_gat), .Y(G7276_1247_ngat) );
INVXL U_g4203 (.A(G7279_1595_gat), .Y(G7279_1595_ngat) );
INVXL U_g4204 (.A(G7420_1249_gat), .Y(G7420_1249_ngat) );
INVXL U_g4205 (.A(G7423_1687_gat), .Y(G7423_1687_ngat) );
INVXL U_g4206 (.A(G6792_1252_gat), .Y(G6792_1252_ngat) );
INVXL U_g4207 (.A(G6795_1591_gat), .Y(G6795_1591_ngat) );
INVXL U_g4208 (.A(G6789_1253_gat), .Y(G6789_1253_ngat) );
INVXL U_g4209 (.A(G6796_1590_gat), .Y(G6796_1590_ngat) );
INVXL U_g4210 (.A(G7380_1257_gat), .Y(G7380_1257_ngat) );
INVXL U_g4211 (.A(G7383_1685_gat), .Y(G7383_1685_ngat) );
INVXL U_g4212 (.A(G7273_1258_gat), .Y(G7273_1258_ngat) );
INVXL U_g4213 (.A(G7280_1586_gat), .Y(G7280_1586_ngat) );
INVXL U_g4214 (.A(G6802_1261_gat), .Y(G6802_1261_ngat) );
INVXL U_g4215 (.A(G6805_1624_gat), .Y(G6805_1624_ngat) );
INVXL U_g4216 (.A(G7372_1263_gat), .Y(G7372_1263_ngat) );
INVXL U_g4217 (.A(G7375_1682_gat), .Y(G7375_1682_ngat) );
INVXL U_g4218 (.A(G7286_1264_gat), .Y(G7286_1264_ngat) );
INVXL U_g4219 (.A(G7289_1628_gat), .Y(G7289_1628_ngat) );
INVXL U_g4220 (.A(G6740_1265_gat), .Y(G6740_1265_ngat) );
INVXL U_g4221 (.A(G6743_1693_gat), .Y(G6743_1693_ngat) );
INVXL U_g4222 (.A(G6474_1269_gat), .Y(G6474_1269_ngat) );
INVXL U_g4223 (.A(G6477_1639_gat), .Y(G6477_1639_ngat) );
INVXL U_g4224 (.A(G6506_1272_gat), .Y(G6506_1272_ngat) );
INVXL U_g4225 (.A(G6509_1649_gat), .Y(G6509_1649_ngat) );
INVXL U_g4226 (.A(G7208_978_gat), .Y(G7208_978_ngat) );
INVXL U_g4227 (.A(G7211_1609_gat), .Y(G7211_1609_ngat) );
INVXL U_g4228 (.A(G6724_979_gat), .Y(G6724_979_ngat) );
INVXL U_g4229 (.A(G6727_1611_gat), .Y(G6727_1611_ngat) );
INVXL U_g4230 (.A(G825_1279_gat), .Y(G825_1279_ngat) );
INVXL U_g4231 (.A(G826_1614_gat), .Y(G826_1614_ngat) );
INVXL U_g4232 (.A(G1053_1280_gat), .Y(G1053_1280_ngat) );
INVXL U_g4233 (.A(G1054_1615_gat), .Y(G1054_1615_ngat) );
INVXL U_g4234 (.A(G3193_1731_gat), .Y(G3193_1731_ngat) );
INVXL U_g4235 (.A(G3194_1617_gat), .Y(G3194_1617_ngat) );
INVXL U_g4236 (.A(G7388_1283_gat), .Y(G7388_1283_ngat) );
INVXL U_g4237 (.A(G7391_1662_gat), .Y(G7391_1662_ngat) );
INVXL U_g4238 (.A(G6781_1286_gat), .Y(G6781_1286_ngat) );
INVXL U_g4239 (.A(G6788_1719_gat), .Y(G6788_1719_ngat) );
INVXL U_g4240 (.A(G6799_1289_gat), .Y(G6799_1289_ngat) );
INVXL U_g4241 (.A(G6806_1598_gat), .Y(G6806_1598_ngat) );
INVXL U_g4242 (.A(G7364_1292_gat), .Y(G7364_1292_ngat) );
INVXL U_g4243 (.A(G7367_1681_gat), .Y(G7367_1681_ngat) );
INVXL U_g4244 (.A(G7283_1294_gat), .Y(G7283_1294_ngat) );
INVXL U_g4245 (.A(G7290_1600_gat), .Y(G7290_1600_ngat) );
INVXL U_g4246 (.A(G6732_1295_gat), .Y(G6732_1295_ngat) );
INVXL U_g4247 (.A(G6735_1634_gat), .Y(G6735_1634_ngat) );
INVXL U_g4248 (.A(G6490_1299_gat), .Y(G6490_1299_ngat) );
INVXL U_g4249 (.A(G6493_1647_gat), .Y(G6493_1647_ngat) );
INVXL U_g4250 (.A(G7216_1300_gat), .Y(G7216_1300_ngat) );
INVXL U_g4251 (.A(G7219_1638_gat), .Y(G7219_1638_ngat) );
INVXL U_g4252 (.A(G6729_1301_gat), .Y(G6729_1301_ngat) );
INVXL U_g4253 (.A(G6736_1629_gat), .Y(G6736_1629_ngat) );
INVXL U_g4254 (.A(G6482_1304_gat), .Y(G6482_1304_ngat) );
INVXL U_g4255 (.A(G6485_1678_gat), .Y(G6485_1678_ngat) );
INVXL U_g4256 (.A(G7213_1306_gat), .Y(G7213_1306_ngat) );
INVXL U_g4257 (.A(G7220_1633_gat), .Y(G7220_1633_ngat) );
INVXL U_g4258 (.A(G6471_1307_gat), .Y(G6471_1307_ngat) );
INVXL U_g4259 (.A(G6478_1604_gat), .Y(G6478_1604_ngat) );
INVXL U_g4260 (.A(G7570_1308_gat), .Y(G7570_1308_ngat) );
INVXL U_g4261 (.A(G7573_1643_gat), .Y(G7573_1643_ngat) );
INVXL U_g4262 (.A(G7567_1310_gat), .Y(G7567_1310_ngat) );
INVXL U_g4263 (.A(G7574_1640_gat), .Y(G7574_1640_ngat) );
INVXL U_g4264 (.A(G7578_1312_gat), .Y(G7578_1312_ngat) );
INVXL U_g4265 (.A(G7581_1677_gat), .Y(G7581_1677_ngat) );
INVXL U_g4266 (.A(G6487_1313_gat), .Y(G6487_1313_ngat) );
INVXL U_g4267 (.A(G6494_1632_gat), .Y(G6494_1632_ngat) );
INVXL U_g4268 (.A(G7562_1314_gat), .Y(G7562_1314_ngat) );
INVXL U_g4269 (.A(G7565_1679_gat), .Y(G7565_1679_ngat) );
INVXL U_g4270 (.A(G6503_1315_gat), .Y(G6503_1315_ngat) );
INVXL U_g4271 (.A(G6510_1607_gat), .Y(G6510_1607_ngat) );
INVXL U_g4272 (.A(G7515_1317_gat), .Y(G7515_1317_ngat) );
INVXL U_g4273 (.A(G7522_1660_gat), .Y(G7522_1660_ngat) );
INVXL U_g4274 (.A(G7526_1320_gat), .Y(G7526_1320_ngat) );
INVXL U_g4275 (.A(G7529_1661_gat), .Y(G7529_1661_ngat) );
INVXL U_g4276 (.A(G7518_1322_gat), .Y(G7518_1322_ngat) );
INVXL U_g4277 (.A(G7521_1652_gat), .Y(G7521_1652_ngat) );
INVXL U_g4278 (.A(G7523_1323_gat), .Y(G7523_1323_ngat) );
INVXL U_g4279 (.A(G7530_1657_gat), .Y(G7530_1657_ngat) );
INVXL U_g4280 (.A(G7385_1324_gat), .Y(G7385_1324_ngat) );
INVXL U_g4281 (.A(G7392_1618_gat), .Y(G7392_1618_ngat) );
INVXL U_g4282 (.A(G4552_1664_gat), .Y(G4552_1664_ngat) );
INVXL U_g4283 (.A(G4553_1663_gat), .Y(G4553_1663_ngat) );
INVXL U_g4284 (.A(G6755_1328_gat), .Y(G6755_1328_ngat) );
INVXL U_g4285 (.A(G6762_1689_gat), .Y(G6762_1689_ngat) );
INVXL U_g4286 (.A(G7247_1691_gat), .Y(G7247_1691_ngat) );
INVXL U_g4287 (.A(G7248_1668_gat), .Y(G7248_1668_ngat) );
INVXL U_g4288 (.A(G6442_1006_gat), .Y(G6442_1006_ngat) );
INVXL U_g4289 (.A(G6445_1670_gat), .Y(G6445_1670_ngat) );
INVXL U_g4290 (.A(G7585_1334_gat), .Y(G7585_1334_ngat) );
INVXL U_g4291 (.A(G7592_1674_gat), .Y(G7592_1674_ngat) );
INVXL U_g4292 (.A(G7588_1336_gat), .Y(G7588_1336_ngat) );
INVXL U_g4293 (.A(G7591_1671_gat), .Y(G7591_1671_ngat) );
INVXL U_g4294 (.A(G7575_1338_gat), .Y(G7575_1338_ngat) );
INVXL U_g4295 (.A(G7582_1646_gat), .Y(G7582_1646_ngat) );
INVXL U_g4296 (.A(G6479_1339_gat), .Y(G6479_1339_ngat) );
INVXL U_g4297 (.A(G6486_1637_gat), .Y(G6486_1637_ngat) );
INVXL U_g4298 (.A(G7559_1340_gat), .Y(G7559_1340_ngat) );
INVXL U_g4299 (.A(G7566_1648_gat), .Y(G7566_1648_ngat) );
INVXL U_g4300 (.A(G7554_1011_gat), .Y(G7554_1011_ngat) );
INVXL U_g4301 (.A(G7557_1651_gat), .Y(G7557_1651_ngat) );
INVXL U_g4302 (.A(G7541_1342_gat), .Y(G7541_1342_ngat) );
INVXL U_g4303 (.A(G7548_1683_gat), .Y(G7548_1683_ngat) );
INVXL U_g4304 (.A(G7361_1343_gat), .Y(G7361_1343_ngat) );
INVXL U_g4305 (.A(G7368_1627_gat), .Y(G7368_1627_ngat) );
INVXL U_g4306 (.A(G7369_1344_gat), .Y(G7369_1344_ngat) );
INVXL U_g4307 (.A(G7376_1599_gat), .Y(G7376_1599_ngat) );
INVXL U_g4308 (.A(G7544_1345_gat), .Y(G7544_1345_ngat) );
INVXL U_g4309 (.A(G7547_1680_gat), .Y(G7547_1680_ngat) );
INVXL U_g4310 (.A(G7531_1346_gat), .Y(G7531_1346_ngat) );
INVXL U_g4311 (.A(G7538_1686_gat), .Y(G7538_1686_ngat) );
INVXL U_g4312 (.A(G7377_1347_gat), .Y(G7377_1347_ngat) );
INVXL U_g4313 (.A(G7384_1594_gat), .Y(G7384_1594_ngat) );
INVXL U_g4314 (.A(G7534_1348_gat), .Y(G7534_1348_ngat) );
INVXL U_g4315 (.A(G7537_1684_gat), .Y(G7537_1684_ngat) );
INVXL U_g4316 (.A(G7417_1349_gat), .Y(G7417_1349_ngat) );
INVXL U_g4317 (.A(G7424_1587_gat), .Y(G7424_1587_ngat) );
INVXL U_g4318 (.A(G6758_1351_gat), .Y(G6758_1351_ngat) );
INVXL U_g4319 (.A(G6761_1666_gat), .Y(G6761_1666_ngat) );
INVXL U_g4320 (.A(G6450_1017_gat), .Y(G6450_1017_ngat) );
INVXL U_g4321 (.A(G6453_1673_gat), .Y(G6453_1673_ngat) );
INVXL U_g4322 (.A(G6466_1019_gat), .Y(G6466_1019_ngat) );
INVXL U_g4323 (.A(G6469_1642_gat), .Y(G6469_1642_ngat) );
INVXL U_g4324 (.A(G7221_1020_gat), .Y(G7221_1020_ngat) );
INVXL U_g4325 (.A(G7228_1606_gat), .Y(G7228_1606_ngat) );
INVXL U_g4326 (.A(G6737_1360_gat), .Y(G6737_1360_ngat) );
INVXL U_g4327 (.A(G6744_1601_gat), .Y(G6744_1601_ngat) );
INVXL U_g4328 (.A(G4201_1695_gat), .Y(G4201_1695_ngat) );
INVXL U_g4329 (.A(G4202_1362_gat), .Y(G4202_1362_ngat) );
INVXL U_g4330 (.A(G6768_1023_gat), .Y(G6768_1023_ngat) );
INVXL U_g4331 (.A(G6771_1697_gat), .Y(G6771_1697_ngat) );
INVXL U_g4332 (.A(G4973_1548_gat), .Y(G4973_1548_ngat) );
INVXL U_g4333 (.A(G4976_829_gat), .Y(G4976_829_ngat) );
INVXL U_g4334 (.A(G1156_1368_gat), .Y(G1156_1368_ngat) );
INVXL U_g4335 (.A(G1157_1699_gat), .Y(G1157_1699_ngat) );
INVXL U_g4336 (.A(G1152_1369_gat), .Y(G1152_1369_ngat) );
INVXL U_g4337 (.A(G1153_1700_gat), .Y(G1153_1700_ngat) );
INVXL U_g4338 (.A(G4932_1547_gat), .Y(G4932_1547_ngat) );
INVXL U_g4339 (.A(G4935_722_gat), .Y(G4935_722_ngat) );
INVXL U_g4340 (.A(G6498_1032_gat), .Y(G6498_1032_ngat) );
INVXL U_g4341 (.A(G6501_1645_gat), .Y(G6501_1645_ngat) );
INVXL U_g4342 (.A(G7237_1701_gat), .Y(G7237_1701_ngat) );
INVXL U_g4343 (.A(G7238_1708_gat), .Y(G7238_1708_ngat) );
INVXL U_g4344 (.A(G6748_1373_gat), .Y(G6748_1373_ngat) );
INVXL U_g4345 (.A(G6751_1705_gat), .Y(G6751_1705_ngat) );
INVXL U_g4346 (.A(G6745_1376_gat), .Y(G6745_1376_ngat) );
INVXL U_g4347 (.A(G6752_1702_gat), .Y(G6752_1702_ngat) );
INVXL U_g4348 (.A(G6458_1036_gat), .Y(G6458_1036_ngat) );
INVXL U_g4349 (.A(G6461_1676_gat), .Y(G6461_1676_ngat) );
INVXL U_g4350 (.A(G6776_1384_gat), .Y(G6776_1384_ngat) );
INVXL U_g4351 (.A(G6779_1713_gat), .Y(G6779_1713_ngat) );
INVXL U_g4352 (.A(G7412_1039_gat), .Y(G7412_1039_ngat) );
INVXL U_g4353 (.A(G7415_1659_gat), .Y(G7415_1659_ngat) );
INVXL U_g4354 (.A(G4210_1712_gat), .Y(G4210_1712_ngat) );
INVXL U_g4355 (.A(G4211_1716_gat), .Y(G4211_1716_ngat) );
INVXL U_g4356 (.A(G6773_1388_gat), .Y(G6773_1388_ngat) );
INVXL U_g4357 (.A(G6780_1711_gat), .Y(G6780_1711_ngat) );
INVXL U_g4358 (.A(G7404_1042_gat), .Y(G7404_1042_ngat) );
INVXL U_g4359 (.A(G7407_1654_gat), .Y(G7407_1654_ngat) );
INVXL U_g4360 (.A(G6784_1396_gat), .Y(G6784_1396_ngat) );
INVXL U_g4361 (.A(G6787_1621_gat), .Y(G6787_1621_ngat) );
INVXL U_g4362 (.A(G7396_1045_gat), .Y(G7396_1045_ngat) );
INVXL U_g4363 (.A(G7399_1656_gat), .Y(G7399_1656_ngat) );
INVXL U_g4364 (.A(G7268_1046_gat), .Y(G7268_1046_ngat) );
INVXL U_g4365 (.A(G7271_1620_gat), .Y(G7271_1620_ngat) );
INVXL U_g4366 (.A(G7425_1047_gat), .Y(G7425_1047_ngat) );
INVXL U_g4367 (.A(G7432_1724_gat), .Y(G7432_1724_ngat) );
INVXL U_g4368 (.A(G5932_1726_gat), .Y(G5932_1726_ngat) );
INVXL U_g4369 (.A(G5935_1402_gat), .Y(G5935_1402_ngat) );
INVXL U_g4370 (.A(G6052_1725_gat), .Y(G6052_1725_ngat) );
INVXL U_g4371 (.A(G6055_1403_gat), .Y(G6055_1403_ngat) );
INVXL U_g4372 (.A(G1238_1727_gat), .Y(G1238_1727_ngat) );
INVXL U_g4373 (.A(G1239_1734_gat), .Y(G1239_1734_ngat) );
INVXL U_g4374 (.A(G1256_1728_gat), .Y(G1256_1728_ngat) );
INVXL U_g4375 (.A(G1257_1737_gat), .Y(G1257_1737_ngat) );
INVXL U_g4376 (.A(G1247_1732_gat), .Y(G1247_1732_ngat) );
INVXL U_g4377 (.A(G1248_1730_gat), .Y(G1248_1730_ngat) );
INVXL U_g4378 (.A(G7335_1742_gat), .Y(G7335_1742_ngat) );
INVXL U_g4379 (.A(G7336_1739_gat), .Y(G7336_1739_ngat) );
INVXL U_g4380 (.A(G7325_1746_gat), .Y(G7325_1746_ngat) );
INVXL U_g4381 (.A(G7326_1743_gat), .Y(G7326_1743_ngat) );
INVXL U_g4382 (.A(G5347_1750_gat), .Y(G5347_1750_ngat) );
INVXL U_g4383 (.A(G5348_1749_gat), .Y(G5348_1749_ngat) );
INVXL U_g4384 (.A(G5357_1753_gat), .Y(G5357_1753_ngat) );
INVXL U_g4385 (.A(G5358_1752_gat), .Y(G5358_1752_ngat) );
INVXL U_g4386 (.A(G1233_1754_gat), .Y(G1233_1754_ngat) );
INVXL U_g4387 (.A(G1234_1760_gat), .Y(G1234_1760_ngat) );
INVXL U_g4388 (.A(G1224_1756_gat), .Y(G1224_1756_ngat) );
INVXL U_g4389 (.A(G1225_1755_gat), .Y(G1225_1755_ngat) );
INVXL U_g4390 (.A(G1215_1758_gat), .Y(G1215_1758_ngat) );
INVXL U_g4391 (.A(G1216_1757_gat), .Y(G1216_1757_ngat) );
INVXL U_g4392 (.A(G3227_1925_gat), .Y(G3227_1925_ngat) );
INVXL U_g4393 (.A(G3220_1761_gat), .Y(G3220_1761_ngat) );
INVXL U_g4394 (.A(G3843_1463_gat), .Y(G3843_1463_ngat) );
INVXL U_g4395 (.A(G3844_1762_gat), .Y(G3844_1762_ngat) );
INVXL U_g4396 (.A(G3281_1464_gat), .Y(G3281_1464_ngat) );
INVXL U_g4397 (.A(G3282_1763_gat), .Y(G3282_1763_ngat) );
INVXL U_g4398 (.A(G3293_1465_gat), .Y(G3293_1465_ngat) );
INVXL U_g4399 (.A(G3294_1764_gat), .Y(G3294_1764_ngat) );
INVXL U_g4400 (.A(G3854_1466_gat), .Y(G3854_1466_ngat) );
INVXL U_g4401 (.A(G3855_1765_gat), .Y(G3855_1765_ngat) );
INVXL U_g4402 (.A(G3312_1467_gat), .Y(G3312_1467_ngat) );
INVXL U_g4403 (.A(G3313_1766_gat), .Y(G3313_1766_ngat) );
INVXL U_g4404 (.A(G3872_1468_gat), .Y(G3872_1468_ngat) );
INVXL U_g4405 (.A(G3873_1767_gat), .Y(G3873_1767_ngat) );
INVXL U_g4406 (.A(G3987_1472_gat), .Y(G3987_1472_ngat) );
INVXL U_g4407 (.A(G3988_1770_gat), .Y(G3988_1770_ngat) );
INVXL U_g4408 (.A(G3342_1473_gat), .Y(G3342_1473_ngat) );
INVXL U_g4409 (.A(G3343_1771_gat), .Y(G3343_1771_ngat) );
INVXL U_g4410 (.A(G3897_1475_gat), .Y(G3897_1475_ngat) );
INVXL U_g4411 (.A(G3898_1772_gat), .Y(G3898_1772_ngat) );
INVXL U_g4412 (.A(G3351_1476_gat), .Y(G3351_1476_ngat) );
INVXL U_g4413 (.A(G3352_1773_gat), .Y(G3352_1773_ngat) );
INVXL U_g4414 (.A(G3363_1477_gat), .Y(G3363_1477_ngat) );
INVXL U_g4415 (.A(G3364_1774_gat), .Y(G3364_1774_ngat) );
INVXL U_g4416 (.A(G3909_1478_gat), .Y(G3909_1478_ngat) );
INVXL U_g4417 (.A(G3910_1775_gat), .Y(G3910_1775_ngat) );
INVXL U_g4418 (.A(G3930_1479_gat), .Y(G3930_1479_ngat) );
INVXL U_g4419 (.A(G3931_1776_gat), .Y(G3931_1776_ngat) );
INVXL U_g4420 (.A(G3379_1480_gat), .Y(G3379_1480_ngat) );
INVXL U_g4421 (.A(G3380_1777_gat), .Y(G3380_1777_ngat) );
INVXL U_g4422 (.A(G3955_1481_gat), .Y(G3955_1481_ngat) );
INVXL U_g4423 (.A(G3956_1778_gat), .Y(G3956_1778_ngat) );
INVXL U_g4424 (.A(G3397_1482_gat), .Y(G3397_1482_ngat) );
INVXL U_g4425 (.A(G3398_1779_gat), .Y(G3398_1779_ngat) );
INVXL U_g4426 (.A(G3415_1484_gat), .Y(G3415_1484_ngat) );
INVXL U_g4427 (.A(G3416_1781_gat), .Y(G3416_1781_ngat) );
INVXL U_g4428 (.A(G3995_1486_gat), .Y(G3995_1486_ngat) );
INVXL U_g4429 (.A(G3996_1782_gat), .Y(G3996_1782_ngat) );
INVXL U_g4430 (.A(G2587_1487_gat), .Y(G2587_1487_ngat) );
INVXL U_g4431 (.A(G2588_1783_gat), .Y(G2588_1783_ngat) );
INVXL U_g4432 (.A(G2341_1488_gat), .Y(G2341_1488_ngat) );
INVXL U_g4433 (.A(G2342_1784_gat), .Y(G2342_1784_ngat) );
INVXL U_g4434 (.A(G2352_1489_gat), .Y(G2352_1489_ngat) );
INVXL U_g4435 (.A(G2353_1785_gat), .Y(G2353_1785_ngat) );
INVXL U_g4436 (.A(G2598_1490_gat), .Y(G2598_1490_ngat) );
INVXL U_g4437 (.A(G2599_1786_gat), .Y(G2599_1786_ngat) );
INVXL U_g4438 (.A(G2616_1491_gat), .Y(G2616_1491_ngat) );
INVXL U_g4439 (.A(G2617_1787_gat), .Y(G2617_1787_ngat) );
INVXL U_g4440 (.A(G2370_1492_gat), .Y(G2370_1492_ngat) );
INVXL U_g4441 (.A(G2371_1788_gat), .Y(G2371_1788_ngat) );
INVXL U_g4442 (.A(G2732_1496_gat), .Y(G2732_1496_ngat) );
INVXL U_g4443 (.A(G2733_1791_gat), .Y(G2733_1791_ngat) );
INVXL U_g4444 (.A(G2398_1497_gat), .Y(G2398_1497_ngat) );
INVXL U_g4445 (.A(G2399_1792_gat), .Y(G2399_1792_ngat) );
INVXL U_g4446 (.A(G2407_1499_gat), .Y(G2407_1499_ngat) );
INVXL U_g4447 (.A(G2408_1793_gat), .Y(G2408_1793_ngat) );
INVXL U_g4448 (.A(G2641_1500_gat), .Y(G2641_1500_ngat) );
INVXL U_g4449 (.A(G2642_1794_gat), .Y(G2642_1794_ngat) );
INVXL U_g4450 (.A(G2653_1501_gat), .Y(G2653_1501_ngat) );
INVXL U_g4451 (.A(G2654_1795_gat), .Y(G2654_1795_ngat) );
INVXL U_g4452 (.A(G2418_1502_gat), .Y(G2418_1502_ngat) );
INVXL U_g4453 (.A(G2419_1796_gat), .Y(G2419_1796_ngat) );
INVXL U_g4454 (.A(G2434_1503_gat), .Y(G2434_1503_ngat) );
INVXL U_g4455 (.A(G2435_1797_gat), .Y(G2435_1797_ngat) );
INVXL U_g4456 (.A(G2674_1504_gat), .Y(G2674_1504_ngat) );
INVXL U_g4457 (.A(G2675_1798_gat), .Y(G2675_1798_ngat) );
INVXL U_g4458 (.A(G2699_1505_gat), .Y(G2699_1505_ngat) );
INVXL U_g4459 (.A(G2700_1799_gat), .Y(G2700_1799_ngat) );
INVXL U_g4460 (.A(G2452_1506_gat), .Y(G2452_1506_ngat) );
INVXL U_g4461 (.A(G2453_1800_gat), .Y(G2453_1800_ngat) );
INVXL U_g4462 (.A(G7281_1860_gat), .Y(G7281_1860_ngat) );
INVXL U_g4463 (.A(G7282_1865_gat), .Y(G7282_1865_ngat) );
INVXL U_g4464 (.A(G4350_1861_gat), .Y(G4350_1861_ngat) );
INVXL U_g4465 (.A(G4351_1917_gat), .Y(G4351_1917_ngat) );
INVXL U_g4466 (.A(G6797_1862_gat), .Y(G6797_1862_ngat) );
INVXL U_g4467 (.A(G6798_1863_gat), .Y(G6798_1863_ngat) );
INVXL U_g4468 (.A(G4306_1864_gat), .Y(G4306_1864_ngat) );
INVXL U_g4469 (.A(G4307_1915_gat), .Y(G4307_1915_ngat) );
INVXL U_g4470 (.A(G6807_1866_gat), .Y(G6807_1866_ngat) );
INVXL U_g4471 (.A(G6808_1879_gat), .Y(G6808_1879_ngat) );
INVXL U_g4472 (.A(G4298_1867_gat), .Y(G4298_1867_ngat) );
INVXL U_g4473 (.A(G4299_1912_gat), .Y(G4299_1912_ngat) );
INVXL U_g4474 (.A(G7291_1868_gat), .Y(G7291_1868_ngat) );
INVXL U_g4475 (.A(G7292_1881_gat), .Y(G7292_1881_ngat) );
INVXL U_g4476 (.A(G3543_1869_gat), .Y(G3543_1869_ngat) );
INVXL U_g4477 (.A(G3544_1922_gat), .Y(G3544_1922_ngat) );
INVXL U_g4478 (.A(G3091_1870_gat), .Y(G3091_1870_ngat) );
INVXL U_g4479 (.A(G3092_1888_gat), .Y(G3092_1888_ngat) );
INVXL U_g4480 (.A(G4196_1605_gat), .Y(G4196_1605_ngat) );
INVXL U_g4481 (.A(G4197_1921_gat), .Y(G4197_1921_ngat) );
INVXL U_g4482 (.A(G3120_1871_gat), .Y(G3120_1871_ngat) );
INVXL U_g4483 (.A(G3121_1894_gat), .Y(G3121_1894_ngat) );
INVXL U_g4484 (.A(G4178_1872_gat), .Y(G4178_1872_ngat) );
INVXL U_g4485 (.A(G4179_1608_gat), .Y(G4179_1608_ngat) );
INVXL U_g4486 (.A(G3525_1873_gat), .Y(G3525_1873_ngat) );
INVXL U_g4487 (.A(G3526_1610_gat), .Y(G3526_1610_ngat) );
INVXL U_g4488 (.A(G4315_1877_gat), .Y(G4315_1877_ngat) );
INVXL U_g4489 (.A(G4316_1899_gat), .Y(G4316_1899_ngat) );
INVXL U_g4490 (.A(G4219_1942_gat), .Y(G4219_1942_ngat) );
INVXL U_g4491 (.A(G4220_1619_gat), .Y(G4220_1619_ngat) );
INVXL U_g4492 (.A(G3566_1940_gat), .Y(G3566_1940_ngat) );
INVXL U_g4493 (.A(G3567_1878_gat), .Y(G3567_1878_ngat) );
INVXL U_g4494 (.A(G4289_1880_gat), .Y(G4289_1880_ngat) );
INVXL U_g4495 (.A(G4290_1911_gat), .Y(G4290_1911_ngat) );
INVXL U_g4496 (.A(G3534_1882_gat), .Y(G3534_1882_ngat) );
INVXL U_g4497 (.A(G3535_1885_gat), .Y(G3535_1885_ngat) );
INVXL U_g4498 (.A(G3108_1883_gat), .Y(G3108_1883_ngat) );
INVXL U_g4499 (.A(G3109_1892_gat), .Y(G3109_1892_ngat) );
INVXL U_g4500 (.A(G4187_1884_gat), .Y(G4187_1884_ngat) );
INVXL U_g4501 (.A(G4188_1887_gat), .Y(G4188_1887_ngat) );
INVXL U_g4502 (.A(G3100_1886_gat), .Y(G3100_1886_ngat) );
INVXL U_g4503 (.A(G3101_1907_gat), .Y(G3101_1907_ngat) );
INVXL U_g4504 (.A(G4593_1889_gat), .Y(G4593_1889_ngat) );
INVXL U_g4505 (.A(G4594_1890_gat), .Y(G4594_1890_ngat) );
INVXL U_g4506 (.A(G3080_1920_gat), .Y(G3080_1920_ngat) );
INVXL U_g4507 (.A(G3081_1641_gat), .Y(G3081_1641_ngat) );
INVXL U_g4508 (.A(G3117_1930_gat), .Y(G3117_1930_ngat) );
INVXL U_g4509 (.A(G3118_1644_gat), .Y(G3118_1644_ngat) );
INVXL U_g4510 (.A(G7583_1891_gat), .Y(G7583_1891_ngat) );
INVXL U_g4511 (.A(G7584_1906_gat), .Y(G7584_1906_ngat) );
INVXL U_g4512 (.A(G4584_1893_gat), .Y(G4584_1893_ngat) );
INVXL U_g4513 (.A(G4585_1908_gat), .Y(G4585_1908_ngat) );
INVXL U_g4514 (.A(G4575_1909_gat), .Y(G4575_1909_ngat) );
INVXL U_g4515 (.A(G4576_1650_gat), .Y(G4576_1650_ngat) );
INVXL U_g4516 (.A(G4561_1897_gat), .Y(G4561_1897_ngat) );
INVXL U_g4517 (.A(G4562_1895_gat), .Y(G4562_1895_ngat) );
INVXL U_g4518 (.A(G4334_1939_gat), .Y(G4334_1939_ngat) );
INVXL U_g4519 (.A(G4335_1653_gat), .Y(G4335_1653_ngat) );
INVXL U_g4520 (.A(G4325_1941_gat), .Y(G4325_1941_ngat) );
INVXL U_g4521 (.A(G4326_1655_gat), .Y(G4326_1655_ngat) );
INVXL U_g4522 (.A(G4570_1896_gat), .Y(G4570_1896_ngat) );
INVXL U_g4523 (.A(G4571_1898_gat), .Y(G4571_1898_ngat) );
INVXL U_g4524 (.A(G4342_1936_gat), .Y(G4342_1936_ngat) );
INVXL U_g4525 (.A(G4343_1658_gat), .Y(G4343_1658_ngat) );
INVXL U_g4526 (.A(G6763_1918_gat), .Y(G6763_1918_ngat) );
INVXL U_g4527 (.A(G6764_1901_gat), .Y(G6764_1901_ngat) );
INVXL U_g4528 (.A(G3050_1903_gat), .Y(G3050_1903_ngat) );
INVXL U_g4529 (.A(G3051_1669_gat), .Y(G3051_1669_ngat) );
INVXL U_g4530 (.A(G7593_1905_gat), .Y(G7593_1905_ngat) );
INVXL U_g4531 (.A(G7594_1904_gat), .Y(G7594_1904_ngat) );
INVXL U_g4532 (.A(G3060_1919_gat), .Y(G3060_1919_ngat) );
INVXL U_g4533 (.A(G3061_1672_gat), .Y(G3061_1672_ngat) );
INVXL U_g4534 (.A(G3069_1934_gat), .Y(G3069_1934_ngat) );
INVXL U_g4535 (.A(G3070_1675_gat), .Y(G3070_1675_ngat) );
INVXL U_g4536 (.A(G7549_1913_gat), .Y(G7549_1913_ngat) );
INVXL U_g4537 (.A(G7550_1910_gat), .Y(G7550_1910_ngat) );
INVXL U_g4538 (.A(G7539_1916_gat), .Y(G7539_1916_ngat) );
INVXL U_g4539 (.A(G7540_1914_gat), .Y(G7540_1914_ngat) );
INVXL U_g4540 (.A(G3548_1924_gat), .Y(G3548_1924_ngat) );
INVXL U_g4541 (.A(G3549_1696_gat), .Y(G3549_1696_ngat) );
INVXL U_g4542 (.A(G4970_718_gat), .Y(G4970_718_ngat) );
INVXL U_g4543 (.A(G4977_1835_gat), .Y(G4977_1835_ngat) );
INVXL U_g4544 (.A(G4929_564_gat), .Y(G4929_564_ngat) );
INVXL U_g4545 (.A(G4936_1834_gat), .Y(G4936_1834_ngat) );
INVXL U_g4546 (.A(G6753_1932_gat), .Y(G6753_1932_ngat) );
INVXL U_g4547 (.A(G6754_1933_gat), .Y(G6754_1933_ngat) );
INVXL U_g4548 (.A(G3557_1935_gat), .Y(G3557_1935_ngat) );
INVXL U_g4549 (.A(G3558_1938_gat), .Y(G3558_1938_ngat) );
INVXL U_g4550 (.A(G4353_1720_gat), .Y(G4353_1720_ngat) );
INVXL U_g4551 (.A(G4354_1943_gat), .Y(G4354_1943_ngat) );
INVXL U_g4552 (.A(G5929_1048_gat), .Y(G5929_1048_ngat) );
INVXL U_g4553 (.A(G5936_1949_gat), .Y(G5936_1949_ngat) );
INVXL U_g4554 (.A(G6049_1049_gat), .Y(G6049_1049_ngat) );
INVXL U_g4555 (.A(G6056_1948_gat), .Y(G6056_1948_ngat) );
INVXL U_g4556 (.A(G7595_1801_gat), .Y(G7595_1801_ngat) );
INVXL U_g4557 (.A(G7602_2021_gat), .Y(G7602_2021_ngat) );
INVXL U_g4558 (.A(G1816_875_gat), .Y(G1816_875_ngat) );
INVXL U_g4559 (.A(G1945_2019_gat), .Y(G1945_2019_ngat) );
INVXL U_g4560 (.A(G1946_2033_gat), .Y(G1946_2033_ngat) );
INVXL U_g4561 (.A(G1567_876_gat), .Y(G1567_876_ngat) );
INVXL U_g4562 (.A(G1712_2014_gat), .Y(G1712_2014_ngat) );
INVXL U_g4563 (.A(G1713_2030_gat), .Y(G1713_2030_ngat) );
INVXL U_g4564 (.A(G1834_878_gat), .Y(G1834_878_ngat) );
INVXL U_g4565 (.A(G1949_2036_gat), .Y(G1949_2036_ngat) );
INVXL U_g4566 (.A(G7598_1809_gat), .Y(G7598_1809_ngat) );
INVXL U_g4567 (.A(G7601_1997_gat), .Y(G7601_1997_ngat) );
INVXL U_g4568 (.A(G5860_2025_gat), .Y(G5860_2025_ngat) );
INVXL U_g4569 (.A(G5863_1520_gat), .Y(G5863_1520_ngat) );
INVXL U_g4570 (.A(G5852_2026_gat), .Y(G5852_2026_ngat) );
INVXL U_g4571 (.A(G5855_1161_gat), .Y(G5855_1161_ngat) );
INVXL U_g4572 (.A(G1624_894_gat), .Y(G1624_894_ngat) );
INVXL U_g4573 (.A(G1737_2056_gat), .Y(G1737_2056_ngat) );
INVXL U_g4574 (.A(G1738_2067_gat), .Y(G1738_2067_ngat) );
INVXL U_g4575 (.A(G1739_2082_gat), .Y(G1739_2082_ngat) );
INVXL U_g4576 (.A(G1647_899_gat), .Y(G1647_899_ngat) );
INVXL U_g4577 (.A(G1743_2070_gat), .Y(G1743_2070_ngat) );
INVXL U_g4578 (.A(G1744_2085_gat), .Y(G1744_2085_ngat) );
INVXL U_g4579 (.A(G821_929_gat), .Y(G821_929_ngat) );
INVXL U_g4580 (.A(G941_2161_gat), .Y(G941_2161_ngat) );
INVXL U_g4581 (.A(G942_2110_gat), .Y(G942_2110_ngat) );
INVXL U_g4582 (.A(G943_2127_gat), .Y(G943_2127_ngat) );
INVXL U_g4583 (.A(G845_980_gat), .Y(G845_980_ngat) );
INVXL U_g4584 (.A(G947_2113_gat), .Y(G947_2113_ngat) );
INVXL U_g4585 (.A(G948_2130_gat), .Y(G948_2130_ngat) );
INVXL U_g4586 (.A(G7337_1902_gat), .Y(G7337_1902_ngat) );
INVXL U_g4587 (.A(G7344_2203_gat), .Y(G7344_2203_ngat) );
INVXL U_g4588 (.A(G4978_1926_gat), .Y(G4978_1926_ngat) );
INVXL U_g4589 (.A(G4979_2200_gat), .Y(G4979_2200_ngat) );
INVXL U_g4590 (.A(G4937_1929_gat), .Y(G4937_1929_ngat) );
INVXL U_g4591 (.A(G4938_2202_gat), .Y(G4938_2202_ngat) );
INVXL U_g4592 (.A(G7340_1931_gat), .Y(G7340_1931_ngat) );
INVXL U_g4593 (.A(G7343_2191_gat), .Y(G7343_2191_ngat) );
INVXL U_g4594 (.A(G2470_1945_gat), .Y(G2470_1945_ngat) );
INVXL U_g4595 (.A(G2471_2209_gat), .Y(G2471_2209_ngat) );
INVXL U_g4596 (.A(G2740_1947_gat), .Y(G2740_1947_ngat) );
INVXL U_g4597 (.A(G2741_2210_gat), .Y(G2741_2210_ngat) );
INVXL U_g4598 (.A(G7353_1954_gat), .Y(G7353_1954_ngat) );
INVXL U_g4599 (.A(G7360_2216_gat), .Y(G7360_2216_ngat) );
INVXL U_g4600 (.A(G7356_1955_gat), .Y(G7356_1955_ngat) );
INVXL U_g4601 (.A(G7359_2215_gat), .Y(G7359_2215_ngat) );
INVXL U_g4602 (.A(G5362_1956_gat), .Y(G5362_1956_ngat) );
INVXL U_g4603 (.A(G5365_2218_gat), .Y(G5365_2218_ngat) );
INVXL U_g4604 (.A(G5359_1957_gat), .Y(G5359_1957_ngat) );
INVXL U_g4605 (.A(G5366_2217_gat), .Y(G5366_2217_ngat) );
INVXL U_g4606 (.A(G3308_1109_gat), .Y(G3308_1109_ngat) );
INVXL U_g4607 (.A(G3441_2240_gat), .Y(G3441_2240_ngat) );
INVXL U_g4608 (.A(G3442_2251_gat), .Y(G3442_2251_ngat) );
INVXL U_g4609 (.A(G3868_1110_gat), .Y(G3868_1110_ngat) );
INVXL U_g4610 (.A(G4014_2241_gat), .Y(G4014_2241_ngat) );
INVXL U_g4611 (.A(G4015_2257_gat), .Y(G4015_2257_ngat) );
INVXL U_g4612 (.A(G3327_1111_gat), .Y(G3327_1111_ngat) );
INVXL U_g4613 (.A(G3445_2254_gat), .Y(G3445_2254_ngat) );
INVXL U_g4614 (.A(G6682_2244_gat), .Y(G6682_2244_ngat) );
INVXL U_g4615 (.A(G6685_1768_gat), .Y(G6685_1768_ngat) );
INVXL U_g4616 (.A(G6674_2245_gat), .Y(G6674_2245_ngat) );
INVXL U_g4617 (.A(G6677_1474_gat), .Y(G6677_1474_ngat) );
INVXL U_g4618 (.A(G3926_1120_gat), .Y(G3926_1120_ngat) );
INVXL U_g4619 (.A(G4039_2275_gat), .Y(G4039_2275_ngat) );
INVXL U_g4620 (.A(G4040_2285_gat), .Y(G4040_2285_ngat) );
INVXL U_g4621 (.A(G4041_2300_gat), .Y(G4041_2300_ngat) );
INVXL U_g4622 (.A(G3949_1122_gat), .Y(G3949_1122_ngat) );
INVXL U_g4623 (.A(G4045_2288_gat), .Y(G4045_2288_ngat) );
INVXL U_g4624 (.A(G4046_2303_gat), .Y(G4046_2303_ngat) );
INVXL U_g4625 (.A(G2366_1130_gat), .Y(G2366_1130_ngat) );
INVXL U_g4626 (.A(G2503_2323_gat), .Y(G2503_2323_ngat) );
INVXL U_g4627 (.A(G2504_2334_gat), .Y(G2504_2334_ngat) );
INVXL U_g4628 (.A(G2612_1131_gat), .Y(G2612_1131_ngat) );
INVXL U_g4629 (.A(G2765_2324_gat), .Y(G2765_2324_ngat) );
INVXL U_g4630 (.A(G2766_2340_gat), .Y(G2766_2340_ngat) );
INVXL U_g4631 (.A(G2384_1132_gat), .Y(G2384_1132_ngat) );
INVXL U_g4632 (.A(G2507_2337_gat), .Y(G2507_2337_ngat) );
INVXL U_g4633 (.A(G5980_2330_gat), .Y(G5980_2330_ngat) );
INVXL U_g4634 (.A(G5983_1789_gat), .Y(G5983_1789_ngat) );
INVXL U_g4635 (.A(G5972_2331_gat), .Y(G5972_2331_ngat) );
INVXL U_g4636 (.A(G5975_1498_gat), .Y(G5975_1498_ngat) );
INVXL U_g4637 (.A(G2670_1141_gat), .Y(G2670_1141_ngat) );
INVXL U_g4638 (.A(G2792_2355_gat), .Y(G2792_2355_ngat) );
INVXL U_g4639 (.A(G2793_2364_gat), .Y(G2793_2364_ngat) );
INVXL U_g4640 (.A(G2794_2528_gat), .Y(G2794_2528_ngat) );
INVXL U_g4641 (.A(G2693_1143_gat), .Y(G2693_1143_ngat) );
INVXL U_g4642 (.A(G2798_2367_gat), .Y(G2798_2367_ngat) );
INVXL U_g4643 (.A(G2799_2531_gat), .Y(G2799_2531_ngat) );
INVXL U_g4644 (.A(G7436_2394_gat), .Y(G7436_2394_ngat) );
INVXL U_g4645 (.A(G7437_2373_gat), .Y(G7437_2373_ngat) );
INVXL U_g4646 (.A(G5817_2384_gat), .Y(G5817_2384_ngat) );
INVXL U_g4647 (.A(G5824_2380_gat), .Y(G5824_2380_ngat) );
INVXL U_g4648 (.A(G5825_2383_gat), .Y(G5825_2383_ngat) );
INVXL U_g4649 (.A(G5832_2381_gat), .Y(G5832_2381_ngat) );
INVXL U_g4650 (.A(G5841_2392_gat), .Y(G5841_2392_ngat) );
INVXL U_g4651 (.A(G5848_2385_gat), .Y(G5848_2385_ngat) );
INVXL U_g4652 (.A(G5833_2393_gat), .Y(G5833_2393_ngat) );
INVXL U_g4653 (.A(G5840_2386_gat), .Y(G5840_2386_ngat) );
INVXL U_g4654 (.A(G5857_1159_gat), .Y(G5857_1159_ngat) );
INVXL U_g4655 (.A(G5864_2397_gat), .Y(G5864_2397_ngat) );
INVXL U_g4656 (.A(G5849_884_gat), .Y(G5849_884_ngat) );
INVXL U_g4657 (.A(G5856_2398_gat), .Y(G5856_2398_ngat) );
INVXL U_g4658 (.A(G5672_2418_gat), .Y(G5672_2418_ngat) );
INVXL U_g4659 (.A(G5675_1541_gat), .Y(G5675_1541_ngat) );
INVXL U_g4660 (.A(G5584_2419_gat), .Y(G5584_2419_ngat) );
INVXL U_g4661 (.A(G5587_1183_gat), .Y(G5587_1183_ngat) );
INVXL U_g4662 (.A(G4980_2511_gat), .Y(G4980_2511_ngat) );
INVXL U_g4663 (.A(G4987_1549_gat), .Y(G4987_1549_ngat) );
INVXL U_g4664 (.A(G4939_2512_gat), .Y(G4939_2512_ngat) );
INVXL U_g4665 (.A(G4946_1837_gat), .Y(G4946_1837_ngat) );
INVXL U_g4666 (.A(G5102_2481_gat), .Y(G5102_2481_ngat) );
INVXL U_g4667 (.A(G5105_1569_gat), .Y(G5105_1569_ngat) );
INVXL U_g4668 (.A(G5014_2482_gat), .Y(G5014_2482_ngat) );
INVXL U_g4669 (.A(G5017_1219_gat), .Y(G5017_1219_ngat) );
INVXL U_g4670 (.A(G7348_2148_gat), .Y(G7348_2148_ngat) );
INVXL U_g4671 (.A(G7351_2471_gat), .Y(G7351_2471_ngat) );
INVXL U_g4672 (.A(G6822_2150_gat), .Y(G6822_2150_ngat) );
INVXL U_g4673 (.A(G6825_2469_gat), .Y(G6825_2469_ngat) );
INVXL U_g4674 (.A(G6819_2152_gat), .Y(G6819_2152_ngat) );
INVXL U_g4675 (.A(G6826_2467_gat), .Y(G6826_2467_ngat) );
INVXL U_g4676 (.A(G7345_2154_gat), .Y(G7345_2154_ngat) );
INVXL U_g4677 (.A(G7352_2464_gat), .Y(G7352_2464_ngat) );
INVXL U_g4678 (.A(G4369_2486_gat), .Y(G4369_2486_ngat) );
INVXL U_g4679 (.A(G89_48_gat), .Y(G89_48_ngat) );
INVXL U_g4680 (.A(G7614_2181_gat), .Y(G7614_2181_ngat) );
INVXL U_g4681 (.A(G7617_2506_gat), .Y(G7617_2506_ngat) );
INVXL U_g4682 (.A(G6809_2190_gat), .Y(G6809_2190_ngat) );
INVXL U_g4683 (.A(G6816_2515_gat), .Y(G6816_2515_ngat) );
INVXL U_g4684 (.A(G6350_2514_gat), .Y(G6350_2514_ngat) );
INVXL U_g4685 (.A(G6351_2505_gat), .Y(G6351_2505_ngat) );
INVXL U_g4686 (.A(G7611_2193_gat), .Y(G7611_2193_ngat) );
INVXL U_g4687 (.A(G7618_2498_gat), .Y(G7618_2498_ngat) );
INVXL U_g4688 (.A(G7603_2196_gat), .Y(G7603_2196_ngat) );
INVXL U_g4689 (.A(G7610_2508_gat), .Y(G7610_2508_ngat) );
INVXL U_g4690 (.A(G7606_2197_gat), .Y(G7606_2197_ngat) );
INVXL U_g4691 (.A(G7609_2507_gat), .Y(G7609_2507_ngat) );
INVXL U_g4692 (.A(G6812_2204_gat), .Y(G6812_2204_ngat) );
INVXL U_g4693 (.A(G6815_2504_gat), .Y(G6815_2504_ngat) );
INVXL U_g4694 (.A(G6340_2539_gat), .Y(G6340_2539_ngat) );
INVXL U_g4695 (.A(G6341_2538_gat), .Y(G6341_2538_ngat) );
INVXL U_g4696 (.A(G5367_2540_gat), .Y(G5367_2540_ngat) );
INVXL U_g4697 (.A(G5368_2541_gat), .Y(G5368_2541_ngat) );
INVXL U_g4698 (.A(G4836_2745_gat), .Y(G4836_2745_ngat) );
INVXL U_g4699 (.A(G4839_316_gat), .Y(G4839_316_ngat) );
INVXL U_g4700 (.A(G2771_2634_gat), .Y(G2771_2634_ngat) );
INVXL U_g4701 (.A(G4526_205_gat), .Y(G4526_205_ngat) );
INVXL U_g4702 (.A(G6639_2560_gat), .Y(G6639_2560_ngat) );
INVXL U_g4703 (.A(G6646_2556_gat), .Y(G6646_2556_ngat) );
INVXL U_g4704 (.A(G6647_2559_gat), .Y(G6647_2559_ngat) );
INVXL U_g4705 (.A(G6654_2557_gat), .Y(G6654_2557_ngat) );
INVXL U_g4706 (.A(G6663_2567_gat), .Y(G6663_2567_ngat) );
INVXL U_g4707 (.A(G6670_2563_gat), .Y(G6670_2563_ngat) );
INVXL U_g4708 (.A(G6655_2568_gat), .Y(G6655_2568_ngat) );
INVXL U_g4709 (.A(G6662_2564_gat), .Y(G6662_2564_ngat) );
INVXL U_g4710 (.A(G6679_1469_gat), .Y(G6679_1469_ngat) );
INVXL U_g4711 (.A(G6686_2570_gat), .Y(G6686_2570_ngat) );
INVXL U_g4712 (.A(G6671_1116_gat), .Y(G6671_1116_ngat) );
INVXL U_g4713 (.A(G6678_2571_gat), .Y(G6678_2571_ngat) );
INVXL U_g4714 (.A(G7132_2589_gat), .Y(G7132_2589_ngat) );
INVXL U_g4715 (.A(G7135_1780_gat), .Y(G7135_1780_ngat) );
INVXL U_g4716 (.A(G7044_2590_gat), .Y(G7044_2590_ngat) );
INVXL U_g4717 (.A(G7047_1485_gat), .Y(G7047_1485_ngat) );
INVXL U_g4718 (.A(G5937_2610_gat), .Y(G5937_2610_ngat) );
INVXL U_g4719 (.A(G5944_2606_gat), .Y(G5944_2606_ngat) );
INVXL U_g4720 (.A(G5945_2609_gat), .Y(G5945_2609_ngat) );
INVXL U_g4721 (.A(G5952_2607_gat), .Y(G5952_2607_ngat) );
INVXL U_g4722 (.A(G5961_2617_gat), .Y(G5961_2617_ngat) );
INVXL U_g4723 (.A(G5968_2613_gat), .Y(G5968_2613_ngat) );
INVXL U_g4724 (.A(G5953_2618_gat), .Y(G5953_2618_ngat) );
INVXL U_g4725 (.A(G5960_2614_gat), .Y(G5960_2614_ngat) );
INVXL U_g4726 (.A(G5977_1493_gat), .Y(G5977_1493_ngat) );
INVXL U_g4727 (.A(G5984_2622_gat), .Y(G5984_2622_ngat) );
INVXL U_g4728 (.A(G5969_1137_gat), .Y(G5969_1137_ngat) );
INVXL U_g4729 (.A(G5976_2623_gat), .Y(G5976_2623_ngat) );
INVXL U_g4730 (.A(G5820_2002_gat), .Y(G5820_2002_ngat) );
INVXL U_g4731 (.A(G5823_2657_gat), .Y(G5823_2657_ngat) );
INVXL U_g4732 (.A(G5828_2003_gat), .Y(G5828_2003_ngat) );
INVXL U_g4733 (.A(G5831_2656_gat), .Y(G5831_2656_ngat) );
INVXL U_g4734 (.A(G5844_2007_gat), .Y(G5844_2007_ngat) );
INVXL U_g4735 (.A(G5847_2663_gat), .Y(G5847_2663_ngat) );
INVXL U_g4736 (.A(G5836_2008_gat), .Y(G5836_2008_ngat) );
INVXL U_g4737 (.A(G5839_2664_gat), .Y(G5839_2664_ngat) );
INVXL U_g4738 (.A(G5526_2662_gat), .Y(G5526_2662_ngat) );
INVXL U_g4739 (.A(G5529_1519_gat), .Y(G5529_1519_ngat) );
INVXL U_g4740 (.A(G2003_2399_gat), .Y(G2003_2399_ngat) );
INVXL U_g4741 (.A(G2004_2666_gat), .Y(G2004_2666_ngat) );
INVXL U_g4742 (.A(G1999_2400_gat), .Y(G1999_2400_ngat) );
INVXL U_g4743 (.A(G2000_2667_gat), .Y(G2000_2667_ngat) );
INVXL U_g4744 (.A(G5468_2665_gat), .Y(G5468_2665_ngat) );
INVXL U_g4745 (.A(G5471_1162_gat), .Y(G5471_1162_ngat) );
INVXL U_g4746 (.A(G4625_2678_gat), .Y(G4625_2678_ngat) );
INVXL U_g4747 (.A(G4626_2404_gat), .Y(G4626_2404_ngat) );
INVXL U_g4748 (.A(G4622_2673_gat), .Y(G4622_2673_ngat) );
INVXL U_g4749 (.A(G4623_2420_gat), .Y(G4623_2420_ngat) );
INVXL U_g4750 (.A(G5669_1182_gat), .Y(G5669_1182_ngat) );
INVXL U_g4751 (.A(G5676_2671_gat), .Y(G5676_2671_ngat) );
INVXL U_g4752 (.A(G5581_911_gat), .Y(G5581_911_ngat) );
INVXL U_g4753 (.A(G5588_2672_gat), .Y(G5588_2672_ngat) );
INVXL U_g4754 (.A(G4983_1191_gat), .Y(G4983_1191_ngat) );
INVXL U_g4755 (.A(G4986_2742_gat), .Y(G4986_2742_ngat) );
INVXL U_g4756 (.A(G4942_1551_gat), .Y(G4942_1551_ngat) );
INVXL U_g4757 (.A(G4945_2743_gat), .Y(G4945_2743_ngat) );
INVXL U_g4758 (.A(G3598_2692_gat), .Y(G3598_2692_ngat) );
INVXL U_g4759 (.A(G3599_2436_gat), .Y(G3599_2436_ngat) );
INVXL U_g4760 (.A(G3595_2688_gat), .Y(G3595_2688_ngat) );
INVXL U_g4761 (.A(G3596_2450_gat), .Y(G3596_2450_ngat) );
INVXL U_g4762 (.A(G5099_1218_gat), .Y(G5099_1218_ngat) );
INVXL U_g4763 (.A(G5106_2712_gat), .Y(G5106_2712_ngat) );
INVXL U_g4764 (.A(G5011_941_gat), .Y(G5011_941_ngat) );
INVXL U_g4765 (.A(G5018_2713_gat), .Y(G5018_2713_ngat) );
INVXL U_g4766 (.A(G4283_2694_gat), .Y(G4283_2694_ngat) );
INVXL U_g4767 (.A(G4284_2456_gat), .Y(G4284_2456_ngat) );
INVXL U_g4768 (.A(G4286_2693_gat), .Y(G4286_2693_ngat) );
INVXL U_g4769 (.A(G4287_2457_gat), .Y(G4287_2457_ngat) );
INVXL U_g4770 (.A(G1320_2696_gat), .Y(G1320_2696_ngat) );
INVXL U_g4771 (.A(G1321_2460_gat), .Y(G1321_2460_ngat) );
INVXL U_g4772 (.A(G1323_2695_gat), .Y(G1323_2695_ngat) );
INVXL U_g4773 (.A(G1324_2461_gat), .Y(G1324_2461_ngat) );
INVXL U_g4774 (.A(G6360_2697_gat), .Y(G6360_2697_ngat) );
INVXL U_g4775 (.A(G6361_2702_gat), .Y(G6361_2702_ngat) );
INVXL U_g4776 (.A(G6827_2700_gat), .Y(G6827_2700_ngat) );
INVXL U_g4777 (.A(G6828_2701_gat), .Y(G6828_2701_ngat) );
INVXL U_g4778 (.A(G7446_2726_gat), .Y(G7446_2726_ngat) );
INVXL U_g4779 (.A(G7447_2735_gat), .Y(G7447_2735_ngat) );
INVXL U_g4780 (.A(G6817_2744_gat), .Y(G6817_2744_ngat) );
INVXL U_g4781 (.A(G6818_2732_gat), .Y(G6818_2732_ngat) );
INVXL U_g4782 (.A(G7456_2737_gat), .Y(G7456_2737_ngat) );
INVXL U_g4783 (.A(G7457_2736_gat), .Y(G7457_2736_ngat) );
INVXL U_g4784 (.A(G6264_2640_gat), .Y(G6264_2640_ngat) );
INVXL U_g4785 (.A(G6267_2208_gat), .Y(G6267_2208_ngat) );
INVXL U_g4786 (.A(G1314_2749_gat), .Y(G1314_2749_ngat) );
INVXL U_g4787 (.A(G1315_2534_gat), .Y(G1315_2534_ngat) );
INVXL U_g4788 (.A(G1317_2748_gat), .Y(G1317_2748_ngat) );
INVXL U_g4789 (.A(G1318_2535_gat), .Y(G1318_2535_ngat) );
INVXL U_g4790 (.A(G1311_2753_gat), .Y(G1311_2753_ngat) );
INVXL U_g4791 (.A(G1312_2542_gat), .Y(G1312_2542_ngat) );
INVXL U_g4792 (.A(G1308_2752_gat), .Y(G1308_2752_ngat) );
INVXL U_g4793 (.A(G1309_2545_gat), .Y(G1309_2545_ngat) );
INVXL U_g4794 (.A(G4833_207_gat), .Y(G4833_207_ngat) );
INVXL U_g4795 (.A(G4840_2879_gat), .Y(G4840_2879_ngat) );
INVXL U_g4796 (.A(G6642_2227_gat), .Y(G6642_2227_ngat) );
INVXL U_g4797 (.A(G6645_2762_gat), .Y(G6645_2762_ngat) );
INVXL U_g4798 (.A(G6650_2228_gat), .Y(G6650_2228_ngat) );
INVXL U_g4799 (.A(G6653_2761_gat), .Y(G6653_2761_ngat) );
INVXL U_g4800 (.A(G6666_2232_gat), .Y(G6666_2232_ngat) );
INVXL U_g4801 (.A(G6669_2767_gat), .Y(G6669_2767_ngat) );
INVXL U_g4802 (.A(G6658_2233_gat), .Y(G6658_2233_ngat) );
INVXL U_g4803 (.A(G6661_2768_gat), .Y(G6661_2768_ngat) );
INVXL U_g4804 (.A(G3487_2574_gat), .Y(G3487_2574_ngat) );
INVXL U_g4805 (.A(G3488_2771_gat), .Y(G3488_2771_ngat) );
INVXL U_g4806 (.A(G6986_2769_gat), .Y(G6986_2769_ngat) );
INVXL U_g4807 (.A(G6989_1769_gat), .Y(G6989_1769_ngat) );
INVXL U_g4808 (.A(G6928_2770_gat), .Y(G6928_2770_ngat) );
INVXL U_g4809 (.A(G6931_1471_gat), .Y(G6931_1471_ngat) );
INVXL U_g4810 (.A(G3483_2577_gat), .Y(G3483_2577_ngat) );
INVXL U_g4811 (.A(G3484_2772_gat), .Y(G3484_2772_ngat) );
INVXL U_g4812 (.A(G7129_1483_gat), .Y(G7129_1483_ngat) );
INVXL U_g4813 (.A(G7136_2776_gat), .Y(G7136_2776_ngat) );
INVXL U_g4814 (.A(G7041_1127_gat), .Y(G7041_1127_ngat) );
INVXL U_g4815 (.A(G7048_2777_gat), .Y(G7048_2777_ngat) );
INVXL U_g4816 (.A(G2761_2783_gat), .Y(G2761_2783_ngat) );
INVXL U_g4817 (.A(G2753_2603_gat), .Y(G2753_2603_ngat) );
INVXL U_g4818 (.A(G5940_2310_gat), .Y(G5940_2310_ngat) );
INVXL U_g4819 (.A(G5943_2791_gat), .Y(G5943_2791_ngat) );
INVXL U_g4820 (.A(G5948_2311_gat), .Y(G5948_2311_ngat) );
INVXL U_g4821 (.A(G5951_2790_gat), .Y(G5951_2790_ngat) );
INVXL U_g4822 (.A(G2499_2782_gat), .Y(G2499_2782_ngat) );
INVXL U_g4823 (.A(G2491_2608_gat), .Y(G2491_2608_ngat) );
INVXL U_g4824 (.A(G5964_2315_gat), .Y(G5964_2315_ngat) );
INVXL U_g4825 (.A(G5967_2796_gat), .Y(G5967_2796_ngat) );
INVXL U_g4826 (.A(G5956_2316_gat), .Y(G5956_2316_ngat) );
INVXL U_g4827 (.A(G5959_2797_gat), .Y(G5959_2797_ngat) );
INVXL U_g4828 (.A(G2559_2624_gat), .Y(G2559_2624_ngat) );
INVXL U_g4829 (.A(G2560_2800_gat), .Y(G2560_2800_ngat) );
INVXL U_g4830 (.A(G6118_2798_gat), .Y(G6118_2798_ngat) );
INVXL U_g4831 (.A(G6121_1790_gat), .Y(G6121_1790_ngat) );
INVXL U_g4832 (.A(G6060_2799_gat), .Y(G6060_2799_ngat) );
INVXL U_g4833 (.A(G6063_1495_gat), .Y(G6063_1495_ngat) );
INVXL U_g4834 (.A(G2555_2627_gat), .Y(G2555_2627_ngat) );
INVXL U_g4835 (.A(G2556_2801_gat), .Y(G2556_2801_ngat) );
INVXL U_g4836 (.A(G4841_2804_gat), .Y(G4841_2804_ngat) );
INVXL U_g4837 (.A(G4848_2631_gat), .Y(G4848_2631_ngat) );
INVXL U_g4838 (.A(G4849_2807_gat), .Y(G4849_2807_ngat) );
INVXL U_g4839 (.A(G4856_2639_gat), .Y(G4856_2639_ngat) );
INVXL U_g4840 (.A(G4857_2810_gat), .Y(G4857_2810_ngat) );
INVXL U_g4841 (.A(G4864_2641_gat), .Y(G4864_2641_ngat) );
INVXL U_g4842 (.A(G4865_2877_gat), .Y(G4865_2877_ngat) );
INVXL U_g4843 (.A(G4872_2649_gat), .Y(G4872_2649_ngat) );
INVXL U_g4844 (.A(G1985_2817_gat), .Y(G1985_2817_ngat) );
INVXL U_g4845 (.A(G1986_2653_gat), .Y(G1986_2653_ngat) );
INVXL U_g4846 (.A(G1988_2818_gat), .Y(G1988_2818_ngat) );
INVXL U_g4847 (.A(G1989_2654_gat), .Y(G1989_2654_ngat) );
INVXL U_g4848 (.A(G1995_2819_gat), .Y(G1995_2819_ngat) );
INVXL U_g4849 (.A(G1996_2658_gat), .Y(G1996_2658_ngat) );
INVXL U_g4850 (.A(G1992_2820_gat), .Y(G1992_2820_ngat) );
INVXL U_g4851 (.A(G1993_2659_gat), .Y(G1993_2659_ngat) );
INVXL U_g4852 (.A(G5523_1158_gat), .Y(G5523_1158_ngat) );
INVXL U_g4853 (.A(G5530_2821_gat), .Y(G5530_2821_ngat) );
INVXL U_g4854 (.A(G5465_885_gat), .Y(G5465_885_ngat) );
INVXL U_g4855 (.A(G5472_2822_gat), .Y(G5472_2822_ngat) );
INVXL U_g4856 (.A(G4627_2827_gat), .Y(G4627_2827_ngat) );
INVXL U_g4857 (.A(G4624_2829_gat), .Y(G4624_2829_ngat) );
INVXL U_g4858 (.A(G5677_2676_gat), .Y(G5677_2676_ngat) );
INVXL U_g4859 (.A(G5678_2832_gat), .Y(G5678_2832_ngat) );
INVXL U_g4860 (.A(G5589_2677_gat), .Y(G5589_2677_ngat) );
INVXL U_g4861 (.A(G5590_2833_gat), .Y(G5590_2833_ngat) );
INVXL U_g4862 (.A(G4988_2834_gat), .Y(G4988_2834_ngat) );
INVXL U_g4863 (.A(G4989_2679_gat), .Y(G4989_2679_ngat) );
INVXL U_g4864 (.A(G4947_2836_gat), .Y(G4947_2836_ngat) );
INVXL U_g4865 (.A(G4948_2680_gat), .Y(G4948_2680_ngat) );
INVXL U_g4866 (.A(G3600_2838_gat), .Y(G3600_2838_ngat) );
INVXL U_g4867 (.A(G3597_2841_gat), .Y(G3597_2841_ngat) );
INVXL U_g4868 (.A(G5107_2690_gat), .Y(G5107_2690_ngat) );
INVXL U_g4869 (.A(G5108_2843_gat), .Y(G5108_2843_ngat) );
INVXL U_g4870 (.A(G5019_2691_gat), .Y(G5019_2691_ngat) );
INVXL U_g4871 (.A(G5020_2844_gat), .Y(G5020_2844_ngat) );
INVXL U_g4872 (.A(G4288_2846_gat), .Y(G4288_2846_ngat) );
INVXL U_g4873 (.A(G4285_2845_gat), .Y(G4285_2845_ngat) );
INVXL U_g4874 (.A(G1325_2848_gat), .Y(G1325_2848_ngat) );
INVXL U_g4875 (.A(G1322_2847_gat), .Y(G1322_2847_ngat) );
INVXL U_g4876 (.A(G4368_2855_gat), .Y(G4368_2855_ngat) );
INVXL U_g4877 (.A(G4360_2699_gat), .Y(G4360_2699_ngat) );
INVXL U_g4878 (.A(G3604_2853_gat), .Y(G3604_2853_ngat) );
INVXL U_g4879 (.A(G3605_2703_gat), .Y(G3605_2703_ngat) );
INVXL U_g4880 (.A(G4274_2852_gat), .Y(G4274_2852_ngat) );
INVXL U_g4881 (.A(G4275_2707_gat), .Y(G4275_2707_ngat) );
INVXL U_g4882 (.A(G4271_2857_gat), .Y(G4271_2857_ngat) );
INVXL U_g4883 (.A(G4272_2710_gat), .Y(G4272_2710_ngat) );
INVXL U_g4884 (.A(G3601_2856_gat), .Y(G3601_2856_ngat) );
INVXL U_g4885 (.A(G3602_2711_gat), .Y(G3602_2711_ngat) );
INVXL U_g4886 (.A(G3610_2873_gat), .Y(G3610_2873_ngat) );
INVXL U_g4887 (.A(G3611_2718_gat), .Y(G3611_2718_ngat) );
INVXL U_g4888 (.A(G4637_2864_gat), .Y(G4637_2864_ngat) );
INVXL U_g4889 (.A(G4638_2723_gat), .Y(G4638_2723_ngat) );
INVXL U_g4890 (.A(G3135_2868_gat), .Y(G3135_2868_ngat) );
INVXL U_g4891 (.A(G3127_2725_gat), .Y(G3127_2725_ngat) );
INVXL U_g4892 (.A(G4634_2863_gat), .Y(G4634_2863_ngat) );
INVXL U_g4893 (.A(G4635_2727_gat), .Y(G4635_2727_ngat) );
INVXL U_g4894 (.A(G4628_2865_gat), .Y(G4628_2865_ngat) );
INVXL U_g4895 (.A(G4629_2730_gat), .Y(G4629_2730_ngat) );
INVXL U_g4896 (.A(G4631_2866_gat), .Y(G4631_2866_ngat) );
INVXL U_g4897 (.A(G4632_2731_gat), .Y(G4632_2731_ngat) );
INVXL U_g4898 (.A(G4277_2876_gat), .Y(G4277_2876_ngat) );
INVXL U_g4899 (.A(G4278_2739_gat), .Y(G4278_2739_ngat) );
INVXL U_g4900 (.A(G4280_2872_gat), .Y(G4280_2872_ngat) );
INVXL U_g4901 (.A(G4281_2740_gat), .Y(G4281_2740_ngat) );
INVXL U_g4902 (.A(G3607_2875_gat), .Y(G3607_2875_ngat) );
INVXL U_g4903 (.A(G3608_2741_gat), .Y(G3608_2741_ngat) );
INVXL U_g4904 (.A(G6261_1944_gat), .Y(G6261_1944_ngat) );
INVXL U_g4905 (.A(G6268_2808_gat), .Y(G6268_2808_ngat) );
INVXL U_g4906 (.A(G6176_2809_gat), .Y(G6176_2809_ngat) );
INVXL U_g4907 (.A(G6179_1946_gat), .Y(G6179_1946_ngat) );
INVXL U_g4908 (.A(G1319_2883_gat), .Y(G1319_2883_ngat) );
INVXL U_g4909 (.A(G1316_2882_gat), .Y(G1316_2882_ngat) );
INVXL U_g4910 (.A(G1313_2886_gat), .Y(G1313_2886_ngat) );
INVXL U_g4911 (.A(G1310_2887_gat), .Y(G1310_2887_ngat) );
INVXL U_g4912 (.A(G3469_2900_gat), .Y(G3469_2900_ngat) );
INVXL U_g4913 (.A(G3470_2758_gat), .Y(G3470_2758_ngat) );
INVXL U_g4914 (.A(G3472_2901_gat), .Y(G3472_2901_ngat) );
INVXL U_g4915 (.A(G3473_2759_gat), .Y(G3473_2759_ngat) );
INVXL U_g4916 (.A(G3479_2902_gat), .Y(G3479_2902_ngat) );
INVXL U_g4917 (.A(G3480_2765_gat), .Y(G3480_2765_ngat) );
INVXL U_g4918 (.A(G3476_2903_gat), .Y(G3476_2903_ngat) );
INVXL U_g4919 (.A(G3477_2766_gat), .Y(G3477_2766_ngat) );
INVXL U_g4920 (.A(G6983_1470_gat), .Y(G6983_1470_ngat) );
INVXL U_g4921 (.A(G6990_2904_gat), .Y(G6990_2904_ngat) );
INVXL U_g4922 (.A(G6925_1115_gat), .Y(G6925_1115_ngat) );
INVXL U_g4923 (.A(G6932_2905_gat), .Y(G6932_2905_ngat) );
INVXL U_g4924 (.A(G7137_2780_gat), .Y(G7137_2780_ngat) );
INVXL U_g4925 (.A(G7138_2913_gat), .Y(G7138_2913_ngat) );
INVXL U_g4926 (.A(G7049_2781_gat), .Y(G7049_2781_ngat) );
INVXL U_g4927 (.A(G7050_2914_gat), .Y(G7050_2914_ngat) );
INVXL U_g4928 (.A(G2541_2918_gat), .Y(G2541_2918_ngat) );
INVXL U_g4929 (.A(G2542_2786_gat), .Y(G2542_2786_ngat) );
INVXL U_g4930 (.A(G2544_2919_gat), .Y(G2544_2919_ngat) );
INVXL U_g4931 (.A(G2545_2787_gat), .Y(G2545_2787_ngat) );
INVXL U_g4932 (.A(G2551_2921_gat), .Y(G2551_2921_ngat) );
INVXL U_g4933 (.A(G2552_2794_gat), .Y(G2552_2794_ngat) );
INVXL U_g4934 (.A(G2548_2922_gat), .Y(G2548_2922_ngat) );
INVXL U_g4935 (.A(G2549_2795_gat), .Y(G2549_2795_ngat) );
INVXL U_g4936 (.A(G6115_1494_gat), .Y(G6115_1494_ngat) );
INVXL U_g4937 (.A(G6122_2923_gat), .Y(G6122_2923_ngat) );
INVXL U_g4938 (.A(G6057_1136_gat), .Y(G6057_1136_ngat) );
INVXL U_g4939 (.A(G6064_2924_gat), .Y(G6064_2924_ngat) );
INVXL U_g4940 (.A(G4844_2345_gat), .Y(G4844_2345_ngat) );
INVXL U_g4941 (.A(G4847_2932_gat), .Y(G4847_2932_ngat) );
INVXL U_g4942 (.A(G4852_2352_gat), .Y(G4852_2352_ngat) );
INVXL U_g4943 (.A(G4855_2935_gat), .Y(G4855_2935_ngat) );
INVXL U_g4944 (.A(G4860_2358_gat), .Y(G4860_2358_ngat) );
INVXL U_g4945 (.A(G4863_2938_gat), .Y(G4863_2938_ngat) );
INVXL U_g4946 (.A(G4868_2371_gat), .Y(G4868_2371_ngat) );
INVXL U_g4947 (.A(G4871_2985_gat), .Y(G4871_2985_ngat) );
INVXL U_g4948 (.A(G7433_2949_gat), .Y(G7433_2949_ngat) );
INVXL U_g4949 (.A(G7442_2814_gat), .Y(G7442_2814_ngat) );
INVXL U_g4950 (.A(G5531_2823_gat), .Y(G5531_2823_ngat) );
INVXL U_g4951 (.A(G5532_2946_gat), .Y(G5532_2946_ngat) );
INVXL U_g4952 (.A(G5473_2826_gat), .Y(G5473_2826_ngat) );
INVXL U_g4953 (.A(G5474_2948_gat), .Y(G5474_2948_ngat) );
INVXL U_g4954 (.A(G5679_2951_gat), .Y(G5679_2951_ngat) );
INVXL U_g4955 (.A(G5686_2830_gat), .Y(G5686_2830_ngat) );
INVXL U_g4956 (.A(G5591_2952_gat), .Y(G5591_2952_ngat) );
INVXL U_g4957 (.A(G5598_2831_gat), .Y(G5598_2831_ngat) );
INVXL U_g4958 (.A(G6829_2957_gat), .Y(G6829_2957_ngat) );
INVXL U_g4959 (.A(G6836_1833_gat), .Y(G6836_1833_ngat) );
INVXL U_g4960 (.A(G4990_2953_gat), .Y(G4990_2953_ngat) );
INVXL U_g4961 (.A(G4997_1555_gat), .Y(G4997_1555_ngat) );
INVXL U_g4962 (.A(G4949_2954_gat), .Y(G4949_2954_ngat) );
INVXL U_g4963 (.A(G4956_1556_gat), .Y(G4956_1556_ngat) );
INVXL U_g4964 (.A(G5109_2959_gat), .Y(G5109_2959_ngat) );
INVXL U_g4965 (.A(G5116_2840_gat), .Y(G5116_2840_ngat) );
INVXL U_g4966 (.A(G5021_2960_gat), .Y(G5021_2960_ngat) );
INVXL U_g4967 (.A(G5028_2842_gat), .Y(G5028_2842_ngat) );
INVXL U_g4968 (.A(G3606_2966_gat), .Y(G3606_2966_ngat) );
INVXL U_g4969 (.A(G3603_2969_gat), .Y(G3603_2969_ngat) );
INVXL U_g4970 (.A(G4276_2967_gat), .Y(G4276_2967_ngat) );
INVXL U_g4971 (.A(G4273_2968_gat), .Y(G4273_2968_ngat) );
INVXL U_g4972 (.A(G3612_2970_gat), .Y(G3612_2970_ngat) );
INVXL U_g4973 (.A(G3609_2984_gat), .Y(G3609_2984_ngat) );
INVXL U_g4974 (.A(G4639_2973_gat), .Y(G4639_2973_ngat) );
INVXL U_g4975 (.A(G4636_2976_gat), .Y(G4636_2976_ngat) );
INVXL U_g4976 (.A(G4633_2978_gat), .Y(G4633_2978_ngat) );
INVXL U_g4977 (.A(G4630_2977_gat), .Y(G4630_2977_ngat) );
INVXL U_g4978 (.A(G4282_2983_gat), .Y(G4282_2983_ngat) );
INVXL U_g4979 (.A(G4279_2982_gat), .Y(G4279_2982_ngat) );
INVXL U_g4980 (.A(G6269_2878_gat), .Y(G6269_2878_ngat) );
INVXL U_g4981 (.A(G6270_2986_gat), .Y(G6270_2986_ngat) );
INVXL U_g4982 (.A(G6173_1723_gat), .Y(G6173_1723_ngat) );
INVXL U_g4983 (.A(G6180_2936_gat), .Y(G6180_2936_ngat) );
INVXL U_g4984 (.A(G5377_2988_gat), .Y(G5377_2988_ngat) );
INVXL U_g4985 (.A(G5384_1953_gat), .Y(G5384_1953_ngat) );
INVXL U_g4986 (.A(G6337_2961_gat), .Y(G6337_2961_ngat) );
INVXL U_g4987 (.A(G6346_2884_gat), .Y(G6346_2884_ngat) );
INVXL U_g4988 (.A(G5385_2962_gat), .Y(G5385_2962_ngat) );
INVXL U_g4989 (.A(G5392_2885_gat), .Y(G5392_2885_ngat) );
INVXL U_g4990 (.A(G5369_2989_gat), .Y(G5369_2989_ngat) );
INVXL U_g4991 (.A(G5376_1961_gat), .Y(G5376_1961_ngat) );
INVXL U_g4992 (.A(G6991_2907_gat), .Y(G6991_2907_ngat) );
INVXL U_g4993 (.A(G6992_3002_gat), .Y(G6992_3002_ngat) );
INVXL U_g4994 (.A(G6933_2908_gat), .Y(G6933_2908_ngat) );
INVXL U_g4995 (.A(G6934_3003_gat), .Y(G6934_3003_ngat) );
INVXL U_g4996 (.A(G7139_3006_gat), .Y(G7139_3006_ngat) );
INVXL U_g4997 (.A(G7146_2911_gat), .Y(G7146_2911_ngat) );
INVXL U_g4998 (.A(G7051_3007_gat), .Y(G7051_3007_ngat) );
INVXL U_g4999 (.A(G7058_2912_gat), .Y(G7058_2912_ngat) );
INVXL U_g5000 (.A(G6123_2926_gat), .Y(G6123_2926_ngat) );
INVXL U_g5001 (.A(G6124_3014_gat), .Y(G6124_3014_ngat) );
INVXL U_g5002 (.A(G6065_2927_gat), .Y(G6065_2927_ngat) );
INVXL U_g5003 (.A(G6066_3015_gat), .Y(G6066_3015_ngat) );
INVXL U_g5004 (.A(G6271_3064_gat), .Y(G6271_3064_ngat) );
INVXL U_g5005 (.A(G6278_2940_gat), .Y(G6278_2940_ngat) );
INVXL U_g5006 (.A(G7438_2650_gat), .Y(G7438_2650_ngat) );
INVXL U_g5007 (.A(G7441_3039_gat), .Y(G7441_3039_ngat) );
INVXL U_g5008 (.A(G5533_3037_gat), .Y(G5533_3037_ngat) );
INVXL U_g5009 (.A(G5540_2660_gat), .Y(G5540_2660_ngat) );
INVXL U_g5010 (.A(G5475_3038_gat), .Y(G5475_3038_ngat) );
INVXL U_g5011 (.A(G5482_2661_gat), .Y(G5482_2661_ngat) );
INVXL U_g5012 (.A(G5682_2674_gat), .Y(G5682_2674_ngat) );
INVXL U_g5013 (.A(G5685_3042_gat), .Y(G5685_3042_ngat) );
INVXL U_g5014 (.A(G5594_2675_gat), .Y(G5594_2675_ngat) );
INVXL U_g5015 (.A(G5597_3043_gat), .Y(G5597_3043_ngat) );
INVXL U_g5016 (.A(G6832_1546_gat), .Y(G6832_1546_ngat) );
INVXL U_g5017 (.A(G6835_3049_gat), .Y(G6835_3049_ngat) );
INVXL U_g5018 (.A(G4993_1203_gat), .Y(G4993_1203_ngat) );
INVXL U_g5019 (.A(G4996_3045_gat), .Y(G4996_3045_ngat) );
INVXL U_g5020 (.A(G4952_1204_gat), .Y(G4952_1204_ngat) );
INVXL U_g5021 (.A(G4955_3046_gat), .Y(G4955_3046_ngat) );
INVXL U_g5022 (.A(G5112_2687_gat), .Y(G5112_2687_ngat) );
INVXL U_g5023 (.A(G5115_3052_gat), .Y(G5115_3052_ngat) );
INVXL U_g5024 (.A(G5024_2689_gat), .Y(G5024_2689_ngat) );
INVXL U_g5025 (.A(G5027_3053_gat), .Y(G5027_3053_ngat) );
INVXL U_g5026 (.A(G6357_3063_gat), .Y(G6357_3063_ngat) );
INVXL U_g5027 (.A(G6366_2963_gat), .Y(G6366_2963_ngat) );
INVXL U_g5028 (.A(G6845_3058_gat), .Y(G6845_3058_ngat) );
INVXL U_g5029 (.A(G6852_2965_gat), .Y(G6852_2965_ngat) );
INVXL U_g5030 (.A(G7443_3061_gat), .Y(G7443_3061_ngat) );
INVXL U_g5031 (.A(G7452_2975_gat), .Y(G7452_2975_ngat) );
INVXL U_g5032 (.A(G6837_3056_gat), .Y(G6837_3056_ngat) );
INVXL U_g5033 (.A(G6844_2979_gat), .Y(G6844_2979_ngat) );
INVXL U_g5034 (.A(G6347_3057_gat), .Y(G6347_3057_ngat) );
INVXL U_g5035 (.A(G6356_2869_gat), .Y(G6356_2869_ngat) );
INVXL U_g5036 (.A(G7453_3062_gat), .Y(G7453_3062_ngat) );
INVXL U_g5037 (.A(G7462_2981_gat), .Y(G7462_2981_ngat) );
INVXL U_g5038 (.A(G6181_2987_gat), .Y(G6181_2987_ngat) );
INVXL U_g5039 (.A(G6182_3065_gat), .Y(G6182_3065_ngat) );
INVXL U_g5040 (.A(G5380_1736_gat), .Y(G5380_1736_ngat) );
INVXL U_g5041 (.A(G5383_3066_gat), .Y(G5383_3066_ngat) );
INVXL U_g5042 (.A(G6342_2750_gat), .Y(G6342_2750_ngat) );
INVXL U_g5043 (.A(G6345_3054_gat), .Y(G6345_3054_ngat) );
INVXL U_g5044 (.A(G5388_2751_gat), .Y(G5388_2751_ngat) );
INVXL U_g5045 (.A(G5391_3055_gat), .Y(G5391_3055_ngat) );
INVXL U_g5046 (.A(G5372_1759_gat), .Y(G5372_1759_ngat) );
INVXL U_g5047 (.A(G5375_3070_gat), .Y(G5375_3070_ngat) );
INVXL U_g5048 (.A(G6993_3076_gat), .Y(G6993_3076_ngat) );
INVXL U_g5049 (.A(G7000_2763_gat), .Y(G7000_2763_ngat) );
INVXL U_g5050 (.A(G6935_3077_gat), .Y(G6935_3077_ngat) );
INVXL U_g5051 (.A(G6942_2764_gat), .Y(G6942_2764_ngat) );
INVXL U_g5052 (.A(G7142_2778_gat), .Y(G7142_2778_ngat) );
INVXL U_g5053 (.A(G7145_3080_gat), .Y(G7145_3080_ngat) );
INVXL U_g5054 (.A(G7054_2779_gat), .Y(G7054_2779_ngat) );
INVXL U_g5055 (.A(G7057_3081_gat), .Y(G7057_3081_ngat) );
INVXL U_g5056 (.A(G6125_3087_gat), .Y(G6125_3087_ngat) );
INVXL U_g5057 (.A(G6132_2792_gat), .Y(G6132_2792_ngat) );
INVXL U_g5058 (.A(G6067_3088_gat), .Y(G6067_3088_ngat) );
INVXL U_g5059 (.A(G6074_2793_gat), .Y(G6074_2793_ngat) );
INVXL U_g5060 (.A(G6183_3131_gat), .Y(G6183_3131_ngat) );
INVXL U_g5061 (.A(G6190_2939_gat), .Y(G6190_2939_ngat) );
INVXL U_g5062 (.A(G6274_2812_gat), .Y(G6274_2812_ngat) );
INVXL U_g5063 (.A(G6277_3130_gat), .Y(G6277_3130_ngat) );
INVXL U_g5064 (.A(G4515_3099_gat), .Y(G4515_3099_ngat) );
INVXL U_g5065 (.A(G4516_3024_gat), .Y(G4516_3024_ngat) );
INVXL U_g5066 (.A(G5536_2387_gat), .Y(G5536_2387_ngat) );
INVXL U_g5067 (.A(G5539_3104_gat), .Y(G5539_3104_ngat) );
INVXL U_g5068 (.A(G5478_2388_gat), .Y(G5478_2388_ngat) );
INVXL U_g5069 (.A(G5481_3105_gat), .Y(G5481_3105_ngat) );
INVXL U_g5070 (.A(G5687_3106_gat), .Y(G5687_3106_ngat) );
INVXL U_g5071 (.A(G5688_3040_gat), .Y(G5688_3040_ngat) );
INVXL U_g5072 (.A(G5599_3107_gat), .Y(G5599_3107_ngat) );
INVXL U_g5073 (.A(G5600_3041_gat), .Y(G5600_3041_ngat) );
INVXL U_g5074 (.A(G3613_3108_gat), .Y(G3613_3108_ngat) );
INVXL U_g5075 (.A(G3614_3044_gat), .Y(G3614_3044_ngat) );
INVXL U_g5076 (.A(G4998_3111_gat), .Y(G4998_3111_ngat) );
INVXL U_g5077 (.A(G4999_3047_gat), .Y(G4999_3047_ngat) );
INVXL U_g5078 (.A(G4957_3112_gat), .Y(G4957_3112_ngat) );
INVXL U_g5079 (.A(G4958_3048_gat), .Y(G4958_3048_ngat) );
INVXL U_g5080 (.A(G3228_2097_gat), .Y(G3228_2097_ngat) );
INVXL U_g5081 (.A(G3242_3098_gat), .Y(G3242_3098_ngat) );
INVXL U_g5082 (.A(G920_2100_gat), .Y(G920_2100_ngat) );
INVXL U_g5083 (.A(G1447_3100_gat), .Y(G1447_3100_ngat) );
INVXL U_g5084 (.A(G5117_3113_gat), .Y(G5117_3113_ngat) );
INVXL U_g5085 (.A(G5118_3050_gat), .Y(G5118_3050_ngat) );
INVXL U_g5086 (.A(G5029_3114_gat), .Y(G5029_3114_ngat) );
INVXL U_g5087 (.A(G5030_3051_gat), .Y(G5030_3051_ngat) );
INVXL U_g5088 (.A(G6362_2849_gat), .Y(G6362_2849_ngat) );
INVXL U_g5089 (.A(G6365_3129_gat), .Y(G6365_3129_ngat) );
INVXL U_g5090 (.A(G6848_2851_gat), .Y(G6848_2851_ngat) );
INVXL U_g5091 (.A(G6851_3120_gat), .Y(G6851_3120_ngat) );
INVXL U_g5092 (.A(G7448_2862_gat), .Y(G7448_2862_ngat) );
INVXL U_g5093 (.A(G7451_3123_gat), .Y(G7451_3123_ngat) );
INVXL U_g5094 (.A(G6840_2867_gat), .Y(G6840_2867_ngat) );
INVXL U_g5095 (.A(G6843_3118_gat), .Y(G6843_3118_ngat) );
INVXL U_g5096 (.A(G6352_2734_gat), .Y(G6352_2734_ngat) );
INVXL U_g5097 (.A(G6355_3119_gat), .Y(G6355_3119_ngat) );
INVXL U_g5098 (.A(G7458_2870_gat), .Y(G7458_2870_ngat) );
INVXL U_g5099 (.A(G7461_3125_gat), .Y(G7461_3125_ngat) );
INVXL U_g5100 (.A(G1329_3132_gat), .Y(G1329_3132_ngat) );
INVXL U_g5101 (.A(G1330_3067_gat), .Y(G1330_3067_ngat) );
INVXL U_g5102 (.A(G2859_3133_gat), .Y(G2859_3133_ngat) );
INVXL U_g5103 (.A(G2860_3068_gat), .Y(G2860_3068_ngat) );
INVXL U_g5104 (.A(G1332_3134_gat), .Y(G1332_3134_ngat) );
INVXL U_g5105 (.A(G1333_3069_gat), .Y(G1333_3069_ngat) );
INVXL U_g5106 (.A(G1326_3135_gat), .Y(G1326_3135_ngat) );
INVXL U_g5107 (.A(G1327_3071_gat), .Y(G1327_3071_ngat) );
INVXL U_g5108 (.A(G6996_2561_gat), .Y(G6996_2561_ngat) );
INVXL U_g5109 (.A(G6999_3140_gat), .Y(G6999_3140_ngat) );
INVXL U_g5110 (.A(G6938_2562_gat), .Y(G6938_2562_ngat) );
INVXL U_g5111 (.A(G6941_3141_gat), .Y(G6941_3141_ngat) );
INVXL U_g5112 (.A(G7147_3142_gat), .Y(G7147_3142_ngat) );
INVXL U_g5113 (.A(G7148_3078_gat), .Y(G7148_3078_ngat) );
INVXL U_g5114 (.A(G7059_3143_gat), .Y(G7059_3143_ngat) );
INVXL U_g5115 (.A(G7060_3079_gat), .Y(G7060_3079_ngat) );
INVXL U_g5116 (.A(G6128_2611_gat), .Y(G6128_2611_ngat) );
INVXL U_g5117 (.A(G6131_3149_gat), .Y(G6131_3149_ngat) );
INVXL U_g5118 (.A(G6070_2612_gat), .Y(G6070_2612_ngat) );
INVXL U_g5119 (.A(G6073_3150_gat), .Y(G6073_3150_ngat) );
INVXL U_g5120 (.A(G6186_2811_gat), .Y(G6186_2811_ngat) );
INVXL U_g5121 (.A(G6189_3187_gat), .Y(G6189_3187_ngat) );
INVXL U_g5122 (.A(G6279_3155_gat), .Y(G6279_3155_ngat) );
INVXL U_g5123 (.A(G6280_3096_gat), .Y(G6280_3096_ngat) );
INVXL U_g5124 (.A(G5541_3159_gat), .Y(G5541_3159_ngat) );
INVXL U_g5125 (.A(G5542_3102_gat), .Y(G5542_3102_ngat) );
INVXL U_g5126 (.A(G5483_3160_gat), .Y(G5483_3160_ngat) );
INVXL U_g5127 (.A(G5484_3103_gat), .Y(G5484_3103_ngat) );
INVXL U_g5128 (.A(G5689_3164_gat), .Y(G5689_3164_ngat) );
INVXL U_g5129 (.A(G5696_2669_gat), .Y(G5696_2669_ngat) );
INVXL U_g5130 (.A(G5601_3166_gat), .Y(G5601_3166_ngat) );
INVXL U_g5131 (.A(G5608_2670_gat), .Y(G5608_2670_ngat) );
INVXL U_g5132 (.A(G4713_3136_gat), .Y(G4713_3136_ngat) );
INVXL U_g5133 (.A(G4720_2430_gat), .Y(G4720_2430_ngat) );
INVXL U_g5134 (.A(G4959_3170_gat), .Y(G4959_3170_ngat) );
INVXL U_g5135 (.A(G4966_1198_gat), .Y(G4966_1198_ngat) );
INVXL U_g5136 (.A(G5000_3169_gat), .Y(G5000_3169_ngat) );
INVXL U_g5137 (.A(G5007_1201_gat), .Y(G5007_1201_ngat) );
INVXL U_g5138 (.A(G5119_3175_gat), .Y(G5119_3175_ngat) );
INVXL U_g5139 (.A(G5126_2685_gat), .Y(G5126_2685_ngat) );
INVXL U_g5140 (.A(G5031_3178_gat), .Y(G5031_3178_ngat) );
INVXL U_g5141 (.A(G5038_2686_gat), .Y(G5038_2686_ngat) );
INVXL U_g5142 (.A(G4753_3158_gat), .Y(G4753_3158_ngat) );
INVXL U_g5143 (.A(G4760_2455_gat), .Y(G4760_2455_ngat) );
INVXL U_g5144 (.A(G2865_3180_gat), .Y(G2865_3180_ngat) );
INVXL U_g5145 (.A(G2866_3115_gat), .Y(G2866_3115_ngat) );
INVXL U_g5146 (.A(G3619_3181_gat), .Y(G3619_3181_ngat) );
INVXL U_g5147 (.A(G3620_3117_gat), .Y(G3620_3117_ngat) );
INVXL U_g5148 (.A(G3136_2475_gat), .Y(G3136_2475_ngat) );
INVXL U_g5149 (.A(G3149_3182_gat), .Y(G3149_3182_ngat) );
INVXL U_g5150 (.A(G4518_3183_gat), .Y(G4518_3183_ngat) );
INVXL U_g5151 (.A(G4519_3124_gat), .Y(G4519_3124_ngat) );
INVXL U_g5152 (.A(G3616_3184_gat), .Y(G3616_3184_ngat) );
INVXL U_g5153 (.A(G3617_3126_gat), .Y(G3617_3126_ngat) );
INVXL U_g5154 (.A(G2862_3185_gat), .Y(G2862_3185_ngat) );
INVXL U_g5155 (.A(G2863_3127_gat), .Y(G2863_3127_ngat) );
INVXL U_g5156 (.A(G4521_3186_gat), .Y(G4521_3186_ngat) );
INVXL U_g5157 (.A(G4522_3128_gat), .Y(G4522_3128_ngat) );
INVXL U_g5158 (.A(G7001_3193_gat), .Y(G7001_3193_ngat) );
INVXL U_g5159 (.A(G7002_3138_gat), .Y(G7002_3138_ngat) );
INVXL U_g5160 (.A(G6943_3194_gat), .Y(G6943_3194_ngat) );
INVXL U_g5161 (.A(G6944_3139_gat), .Y(G6944_3139_ngat) );
INVXL U_g5162 (.A(G7149_3198_gat), .Y(G7149_3198_ngat) );
INVXL U_g5163 (.A(G7156_2774_gat), .Y(G7156_2774_ngat) );
INVXL U_g5164 (.A(G7061_3199_gat), .Y(G7061_3199_ngat) );
INVXL U_g5165 (.A(G7068_2775_gat), .Y(G7068_2775_ngat) );
INVXL U_g5166 (.A(G4793_3203_gat), .Y(G4793_3203_ngat) );
INVXL U_g5167 (.A(G4800_2598_gat), .Y(G4800_2598_ngat) );
INVXL U_g5168 (.A(G6133_3204_gat), .Y(G6133_3204_ngat) );
INVXL U_g5169 (.A(G6134_3146_gat), .Y(G6134_3146_ngat) );
INVXL U_g5170 (.A(G6075_3205_gat), .Y(G6075_3205_ngat) );
INVXL U_g5171 (.A(G6076_3147_gat), .Y(G6076_3147_ngat) );
INVXL U_g5172 (.A(G6281_3209_gat), .Y(G6281_3209_ngat) );
INVXL U_g5173 (.A(G6288_2805_gat), .Y(G6288_2805_ngat) );
INVXL U_g5174 (.A(G6191_3208_gat), .Y(G6191_3208_ngat) );
INVXL U_g5175 (.A(G6192_3154_gat), .Y(G6192_3154_ngat) );
INVXL U_g5176 (.A(G5543_3212_gat), .Y(G5543_3212_ngat) );
INVXL U_g5177 (.A(G5550_2401_gat), .Y(G5550_2401_ngat) );
INVXL U_g5178 (.A(G5485_3213_gat), .Y(G5485_3213_ngat) );
INVXL U_g5179 (.A(G5492_2402_gat), .Y(G5492_2402_ngat) );
INVXL U_g5180 (.A(G4721_3217_gat), .Y(G4721_3217_ngat) );
INVXL U_g5181 (.A(G4728_2412_gat), .Y(G4728_2412_ngat) );
INVXL U_g5182 (.A(G5692_2413_gat), .Y(G5692_2413_ngat) );
INVXL U_g5183 (.A(G5695_3219_gat), .Y(G5695_3219_ngat) );
INVXL U_g5184 (.A(G5604_2414_gat), .Y(G5604_2414_ngat) );
INVXL U_g5185 (.A(G5607_3221_gat), .Y(G5607_3221_ngat) );
INVXL U_g5186 (.A(G4729_3218_gat), .Y(G4729_3218_ngat) );
INVXL U_g5187 (.A(G4736_2415_gat), .Y(G4736_2415_ngat) );
INVXL U_g5188 (.A(G4737_3220_gat), .Y(G4737_3220_ngat) );
INVXL U_g5189 (.A(G4744_2423_gat), .Y(G4744_2423_ngat) );
INVXL U_g5190 (.A(G4745_3222_gat), .Y(G4745_3222_ngat) );
INVXL U_g5191 (.A(G4752_2425_gat), .Y(G4752_2425_ngat) );
INVXL U_g5192 (.A(G4716_2094_gat), .Y(G4716_2094_ngat) );
INVXL U_g5193 (.A(G4719_3192_gat), .Y(G4719_3192_ngat) );
INVXL U_g5194 (.A(G4962_919_gat), .Y(G4962_919_ngat) );
INVXL U_g5195 (.A(G4965_3227_gat), .Y(G4965_3227_ngat) );
INVXL U_g5196 (.A(G5003_920_gat), .Y(G5003_920_ngat) );
INVXL U_g5197 (.A(G5006_3226_gat), .Y(G5006_3226_ngat) );
INVXL U_g5198 (.A(G4761_3233_gat), .Y(G4761_3233_ngat) );
INVXL U_g5199 (.A(G4768_2442_gat), .Y(G4768_2442_ngat) );
INVXL U_g5200 (.A(G5122_2443_gat), .Y(G5122_2443_ngat) );
INVXL U_g5201 (.A(G5125_3234_gat), .Y(G5125_3234_ngat) );
INVXL U_g5202 (.A(G5034_2444_gat), .Y(G5034_2444_ngat) );
INVXL U_g5203 (.A(G5037_3236_gat), .Y(G5037_3236_ngat) );
INVXL U_g5204 (.A(G4769_3242_gat), .Y(G4769_3242_ngat) );
INVXL U_g5205 (.A(G4776_2445_gat), .Y(G4776_2445_ngat) );
INVXL U_g5206 (.A(G4785_3237_gat), .Y(G4785_3237_ngat) );
INVXL U_g5207 (.A(G4792_2449_gat), .Y(G4792_2449_ngat) );
INVXL U_g5208 (.A(G4756_2139_gat), .Y(G4756_2139_ngat) );
INVXL U_g5209 (.A(G4759_3211_gat), .Y(G4759_3211_ngat) );
INVXL U_g5210 (.A(G4777_3235_gat), .Y(G4777_3235_ngat) );
INVXL U_g5211 (.A(G4784_2485_gat), .Y(G4784_2485_ngat) );
INVXL U_g5212 (.A(G7003_3247_gat), .Y(G7003_3247_ngat) );
INVXL U_g5213 (.A(G7010_2575_gat), .Y(G7010_2575_ngat) );
INVXL U_g5214 (.A(G6945_3248_gat), .Y(G6945_3248_ngat) );
INVXL U_g5215 (.A(G6952_2576_gat), .Y(G6952_2576_ngat) );
INVXL U_g5216 (.A(G4801_3250_gat), .Y(G4801_3250_ngat) );
INVXL U_g5217 (.A(G4808_2583_gat), .Y(G4808_2583_ngat) );
INVXL U_g5218 (.A(G7152_2584_gat), .Y(G7152_2584_ngat) );
INVXL U_g5219 (.A(G7155_3255_gat), .Y(G7155_3255_ngat) );
INVXL U_g5220 (.A(G7064_2585_gat), .Y(G7064_2585_ngat) );
INVXL U_g5221 (.A(G7067_3256_gat), .Y(G7067_3256_ngat) );
INVXL U_g5222 (.A(G4809_3253_gat), .Y(G4809_3253_ngat) );
INVXL U_g5223 (.A(G4816_2586_gat), .Y(G4816_2586_ngat) );
INVXL U_g5224 (.A(G4817_3254_gat), .Y(G4817_3254_ngat) );
INVXL U_g5225 (.A(G4824_2593_gat), .Y(G4824_2593_ngat) );
INVXL U_g5226 (.A(G4825_3257_gat), .Y(G4825_3257_ngat) );
INVXL U_g5227 (.A(G4832_2597_gat), .Y(G4832_2597_ngat) );
INVXL U_g5228 (.A(G4796_2304_gat), .Y(G4796_2304_ngat) );
INVXL U_g5229 (.A(G4799_3259_gat), .Y(G4799_3259_ngat) );
INVXL U_g5230 (.A(G6135_3260_gat), .Y(G6135_3260_ngat) );
INVXL U_g5231 (.A(G6142_2625_gat), .Y(G6142_2625_ngat) );
INVXL U_g5232 (.A(G6077_3261_gat), .Y(G6077_3261_ngat) );
INVXL U_g5233 (.A(G6084_2626_gat), .Y(G6084_2626_ngat) );
INVXL U_g5234 (.A(G6284_2635_gat), .Y(G6284_2635_ngat) );
INVXL U_g5235 (.A(G6287_3264_gat), .Y(G6287_3264_ngat) );
INVXL U_g5236 (.A(G6193_3263_gat), .Y(G6193_3263_ngat) );
INVXL U_g5237 (.A(G6200_2933_gat), .Y(G6200_2933_ngat) );
INVXL U_g5238 (.A(G5546_2038_gat), .Y(G5546_2038_ngat) );
INVXL U_g5239 (.A(G5549_3268_gat), .Y(G5549_3268_ngat) );
INVXL U_g5240 (.A(G5488_2039_gat), .Y(G5488_2039_ngat) );
INVXL U_g5241 (.A(G5491_3269_gat), .Y(G5491_3269_ngat) );
INVXL U_g5242 (.A(G4724_2048_gat), .Y(G4724_2048_ngat) );
INVXL U_g5243 (.A(G4727_3278_gat), .Y(G4727_3278_ngat) );
INVXL U_g5244 (.A(G5697_3276_gat), .Y(G5697_3276_ngat) );
INVXL U_g5245 (.A(G5698_3215_gat), .Y(G5698_3215_ngat) );
INVXL U_g5246 (.A(G5609_3277_gat), .Y(G5609_3277_ngat) );
INVXL U_g5247 (.A(G5610_3216_gat), .Y(G5610_3216_ngat) );
INVXL U_g5248 (.A(G4732_2051_gat), .Y(G4732_2051_ngat) );
INVXL U_g5249 (.A(G4735_3280_gat), .Y(G4735_3280_ngat) );
INVXL U_g5250 (.A(G4740_2066_gat), .Y(G4740_2066_ngat) );
INVXL U_g5251 (.A(G4743_3282_gat), .Y(G4743_3282_ngat) );
INVXL U_g5252 (.A(G4748_2075_gat), .Y(G4748_2075_ngat) );
INVXL U_g5253 (.A(G4751_3284_gat), .Y(G4751_3284_ngat) );
INVXL U_g5254 (.A(G4967_3288_gat), .Y(G4967_3288_ngat) );
INVXL U_g5255 (.A(G4968_3224_gat), .Y(G4968_3224_ngat) );
INVXL U_g5256 (.A(G5008_3289_gat), .Y(G5008_3289_ngat) );
INVXL U_g5257 (.A(G5009_3225_gat), .Y(G5009_3225_ngat) );
INVXL U_g5258 (.A(G4764_2102_gat), .Y(G4764_2102_ngat) );
INVXL U_g5259 (.A(G4767_3297_gat), .Y(G4767_3297_ngat) );
INVXL U_g5260 (.A(G5127_3295_gat), .Y(G5127_3295_ngat) );
INVXL U_g5261 (.A(G5128_3231_gat), .Y(G5128_3231_ngat) );
INVXL U_g5262 (.A(G5039_3296_gat), .Y(G5039_3296_ngat) );
INVXL U_g5263 (.A(G5040_3232_gat), .Y(G5040_3232_ngat) );
INVXL U_g5264 (.A(G4772_2105_gat), .Y(G4772_2105_ngat) );
INVXL U_g5265 (.A(G4775_3303_gat), .Y(G4775_3303_ngat) );
INVXL U_g5266 (.A(G4788_2118_gat), .Y(G4788_2118_ngat) );
INVXL U_g5267 (.A(G4791_3301_gat), .Y(G4791_3301_ngat) );
INVXL U_g5268 (.A(G4780_2168_gat), .Y(G4780_2168_ngat) );
INVXL U_g5269 (.A(G4783_3299_gat), .Y(G4783_3299_ngat) );
INVXL U_g5270 (.A(G7006_2259_gat), .Y(G7006_2259_ngat) );
INVXL U_g5271 (.A(G7009_3312_gat), .Y(G7009_3312_ngat) );
INVXL U_g5272 (.A(G6948_2260_gat), .Y(G6948_2260_ngat) );
INVXL U_g5273 (.A(G6951_3313_gat), .Y(G6951_3313_ngat) );
INVXL U_g5274 (.A(G4804_2266_gat), .Y(G4804_2266_ngat) );
INVXL U_g5275 (.A(G4807_3321_gat), .Y(G4807_3321_ngat) );
INVXL U_g5276 (.A(G7157_3322_gat), .Y(G7157_3322_ngat) );
INVXL U_g5277 (.A(G7158_3251_gat), .Y(G7158_3251_ngat) );
INVXL U_g5278 (.A(G7069_3323_gat), .Y(G7069_3323_ngat) );
INVXL U_g5279 (.A(G7070_3252_gat), .Y(G7070_3252_ngat) );
INVXL U_g5280 (.A(G4812_2269_gat), .Y(G4812_2269_ngat) );
INVXL U_g5281 (.A(G4815_3325_gat), .Y(G4815_3325_ngat) );
INVXL U_g5282 (.A(G4820_2281_gat), .Y(G4820_2281_ngat) );
INVXL U_g5283 (.A(G4823_3327_gat), .Y(G4823_3327_ngat) );
INVXL U_g5284 (.A(G4828_2293_gat), .Y(G4828_2293_ngat) );
INVXL U_g5285 (.A(G4831_3329_gat), .Y(G4831_3329_ngat) );
INVXL U_g5286 (.A(G6138_2342_gat), .Y(G6138_2342_ngat) );
INVXL U_g5287 (.A(G6141_3331_gat), .Y(G6141_3331_ngat) );
INVXL U_g5288 (.A(G6080_2343_gat), .Y(G6080_2343_ngat) );
INVXL U_g5289 (.A(G6083_3332_gat), .Y(G6083_3332_ngat) );
INVXL U_g5290 (.A(G6289_3335_gat), .Y(G6289_3335_ngat) );
INVXL U_g5291 (.A(G6290_3262_gat), .Y(G6290_3262_ngat) );
INVXL U_g5292 (.A(G6196_2806_gat), .Y(G6196_2806_ngat) );
INVXL U_g5293 (.A(G6199_3337_gat), .Y(G6199_3337_ngat) );
INVXL U_g5294 (.A(G5551_3344_gat), .Y(G5551_3344_ngat) );
INVXL U_g5295 (.A(G5552_3272_gat), .Y(G5552_3272_ngat) );
INVXL U_g5296 (.A(G5493_3345_gat), .Y(G5493_3345_ngat) );
INVXL U_g5297 (.A(G5494_3273_gat), .Y(G5494_3273_ngat) );
INVXL U_g5298 (.A(G5699_3347_gat), .Y(G5699_3347_ngat) );
INVXL U_g5299 (.A(G5706_2428_gat), .Y(G5706_2428_ngat) );
INVXL U_g5300 (.A(G5611_3348_gat), .Y(G5611_3348_ngat) );
INVXL U_g5301 (.A(G5618_2429_gat), .Y(G5618_2429_ngat) );
INVXL U_g5302 (.A(G5129_3359_gat), .Y(G5129_3359_ngat) );
INVXL U_g5303 (.A(G5136_2453_gat), .Y(G5136_2453_ngat) );
INVXL U_g5304 (.A(G5041_3360_gat), .Y(G5041_3360_ngat) );
INVXL U_g5305 (.A(G5048_2454_gat), .Y(G5048_2454_ngat) );
INVXL U_g5306 (.A(G7011_3373_gat), .Y(G7011_3373_ngat) );
INVXL U_g5307 (.A(G7012_3315_gat), .Y(G7012_3315_ngat) );
INVXL U_g5308 (.A(G6953_3374_gat), .Y(G6953_3374_ngat) );
INVXL U_g5309 (.A(G6954_3316_gat), .Y(G6954_3316_ngat) );
INVXL U_g5310 (.A(G7159_3377_gat), .Y(G7159_3377_ngat) );
INVXL U_g5311 (.A(G7166_2599_gat), .Y(G7166_2599_ngat) );
INVXL U_g5312 (.A(G7071_3378_gat), .Y(G7071_3378_ngat) );
INVXL U_g5313 (.A(G7078_2600_gat), .Y(G7078_2600_ngat) );
INVXL U_g5314 (.A(G6143_3383_gat), .Y(G6143_3383_ngat) );
INVXL U_g5315 (.A(G6144_3333_gat), .Y(G6144_3333_ngat) );
INVXL U_g5316 (.A(G6085_3384_gat), .Y(G6085_3384_ngat) );
INVXL U_g5317 (.A(G6086_3334_gat), .Y(G6086_3334_ngat) );
INVXL U_g5318 (.A(G6201_3386_gat), .Y(G6201_3386_ngat) );
INVXL U_g5319 (.A(G6202_3336_gat), .Y(G6202_3336_ngat) );
INVXL U_g5320 (.A(G5495_3392_gat), .Y(G5495_3392_ngat) );
INVXL U_g5321 (.A(G5502_2395_gat), .Y(G5502_2395_ngat) );
INVXL U_g5322 (.A(G5553_3391_gat), .Y(G5553_3391_ngat) );
INVXL U_g5323 (.A(G5560_2396_gat), .Y(G5560_2396_ngat) );
INVXL U_g5324 (.A(G5702_2090_gat), .Y(G5702_2090_ngat) );
INVXL U_g5325 (.A(G5705_3394_gat), .Y(G5705_3394_ngat) );
INVXL U_g5326 (.A(G5614_2091_gat), .Y(G5614_2091_ngat) );
INVXL U_g5327 (.A(G5617_3395_gat), .Y(G5617_3395_ngat) );
INVXL U_g5328 (.A(G5132_2135_gat), .Y(G5132_2135_ngat) );
INVXL U_g5329 (.A(G5135_3409_gat), .Y(G5135_3409_ngat) );
INVXL U_g5330 (.A(G5044_2136_gat), .Y(G5044_2136_ngat) );
INVXL U_g5331 (.A(G5047_3410_gat), .Y(G5047_3410_ngat) );
INVXL U_g5332 (.A(G6291_3385_gat), .Y(G6291_3385_ngat) );
INVXL U_g5333 (.A(G6298_2880_gat), .Y(G6298_2880_ngat) );
INVXL U_g5334 (.A(G6955_3423_gat), .Y(G6955_3423_ngat) );
INVXL U_g5335 (.A(G6962_2572_gat), .Y(G6962_2572_ngat) );
INVXL U_g5336 (.A(G7013_3422_gat), .Y(G7013_3422_ngat) );
INVXL U_g5337 (.A(G7020_2573_gat), .Y(G7020_2573_ngat) );
INVXL U_g5338 (.A(G7162_2305_gat), .Y(G7162_2305_ngat) );
INVXL U_g5339 (.A(G7165_3427_gat), .Y(G7165_3427_ngat) );
INVXL U_g5340 (.A(G7074_2306_gat), .Y(G7074_2306_ngat) );
INVXL U_g5341 (.A(G7077_3428_gat), .Y(G7077_3428_ngat) );
INVXL U_g5342 (.A(G6087_3435_gat), .Y(G6087_3435_ngat) );
INVXL U_g5343 (.A(G6094_2620_gat), .Y(G6094_2620_ngat) );
INVXL U_g5344 (.A(G6145_3434_gat), .Y(G6145_3434_ngat) );
INVXL U_g5345 (.A(G6152_2621_gat), .Y(G6152_2621_ngat) );
INVXL U_g5346 (.A(G5498_2023_gat), .Y(G5498_2023_ngat) );
INVXL U_g5347 (.A(G5501_3441_gat), .Y(G5501_3441_ngat) );
INVXL U_g5348 (.A(G5556_2024_gat), .Y(G5556_2024_ngat) );
INVXL U_g5349 (.A(G5559_3440_gat), .Y(G5559_3440_ngat) );
INVXL U_g5350 (.A(G5707_3442_gat), .Y(G5707_3442_ngat) );
INVXL U_g5351 (.A(G5708_3399_gat), .Y(G5708_3399_ngat) );
INVXL U_g5352 (.A(G5619_3443_gat), .Y(G5619_3443_ngat) );
INVXL U_g5353 (.A(G5620_3400_gat), .Y(G5620_3400_ngat) );
INVXL U_g5354 (.A(G5137_3447_gat), .Y(G5137_3447_ngat) );
INVXL U_g5355 (.A(G5138_3413_gat), .Y(G5138_3413_ngat) );
INVXL U_g5356 (.A(G5049_3448_gat), .Y(G5049_3448_ngat) );
INVXL U_g5357 (.A(G5050_3414_gat), .Y(G5050_3414_ngat) );
INVXL U_g5358 (.A(G6294_2746_gat), .Y(G6294_2746_ngat) );
INVXL U_g5359 (.A(G6297_3436_gat), .Y(G6297_3436_ngat) );
INVXL U_g5360 (.A(G6203_3437_gat), .Y(G6203_3437_ngat) );
INVXL U_g5361 (.A(G6210_2881_gat), .Y(G6210_2881_ngat) );
INVXL U_g5362 (.A(G6958_2248_gat), .Y(G6958_2248_ngat) );
INVXL U_g5363 (.A(G6961_3457_gat), .Y(G6961_3457_ngat) );
INVXL U_g5364 (.A(G7016_2249_gat), .Y(G7016_2249_ngat) );
INVXL U_g5365 (.A(G7019_3456_gat), .Y(G7019_3456_ngat) );
INVXL U_g5366 (.A(G7167_3458_gat), .Y(G7167_3458_ngat) );
INVXL U_g5367 (.A(G7168_3432_gat), .Y(G7168_3432_ngat) );
INVXL U_g5368 (.A(G7079_3459_gat), .Y(G7079_3459_ngat) );
INVXL U_g5369 (.A(G7080_3433_gat), .Y(G7080_3433_ngat) );
INVXL U_g5370 (.A(G6090_2328_gat), .Y(G6090_2328_ngat) );
INVXL U_g5371 (.A(G6093_3463_gat), .Y(G6093_3463_ngat) );
INVXL U_g5372 (.A(G6148_2329_gat), .Y(G6148_2329_ngat) );
INVXL U_g5373 (.A(G6151_3462_gat), .Y(G6151_3462_ngat) );
INVXL U_g5374 (.A(G5503_3465_gat), .Y(G5503_3465_ngat) );
INVXL U_g5375 (.A(G5504_3438_gat), .Y(G5504_3438_ngat) );
INVXL U_g5376 (.A(G5561_3466_gat), .Y(G5561_3466_ngat) );
INVXL U_g5377 (.A(G5562_3439_gat), .Y(G5562_3439_ngat) );
INVXL U_g5378 (.A(G5621_3468_gat), .Y(G5621_3468_ngat) );
INVXL U_g5379 (.A(G5628_2426_gat), .Y(G5628_2426_ngat) );
INVXL U_g5380 (.A(G5709_3467_gat), .Y(G5709_3467_ngat) );
INVXL U_g5381 (.A(G5716_2427_gat), .Y(G5716_2427_ngat) );
INVXL U_g5382 (.A(G5051_3471_gat), .Y(G5051_3471_ngat) );
INVXL U_g5383 (.A(G5058_2451_gat), .Y(G5058_2451_ngat) );
INVXL U_g5384 (.A(G5139_3470_gat), .Y(G5139_3470_ngat) );
INVXL U_g5385 (.A(G5146_2452_gat), .Y(G5146_2452_ngat) );
INVXL U_g5386 (.A(G6299_3472_gat), .Y(G6299_3472_ngat) );
INVXL U_g5387 (.A(G6300_3453_gat), .Y(G6300_3453_ngat) );
INVXL U_g5388 (.A(G6206_2747_gat), .Y(G6206_2747_ngat) );
INVXL U_g5389 (.A(G6209_3464_gat), .Y(G6209_3464_ngat) );
INVXL U_g5390 (.A(G6963_3474_gat), .Y(G6963_3474_ngat) );
INVXL U_g5391 (.A(G6964_3454_gat), .Y(G6964_3454_ngat) );
INVXL U_g5392 (.A(G7021_3475_gat), .Y(G7021_3475_ngat) );
INVXL U_g5393 (.A(G7022_3455_gat), .Y(G7022_3455_ngat) );
INVXL U_g5394 (.A(G7081_3477_gat), .Y(G7081_3477_ngat) );
INVXL U_g5395 (.A(G7088_2595_gat), .Y(G7088_2595_ngat) );
INVXL U_g5396 (.A(G7169_3476_gat), .Y(G7169_3476_ngat) );
INVXL U_g5397 (.A(G7176_2596_gat), .Y(G7176_2596_ngat) );
INVXL U_g5398 (.A(G6095_3478_gat), .Y(G6095_3478_ngat) );
INVXL U_g5399 (.A(G6096_3460_gat), .Y(G6096_3460_ngat) );
INVXL U_g5400 (.A(G6153_3479_gat), .Y(G6153_3479_ngat) );
INVXL U_g5401 (.A(G6154_3461_gat), .Y(G6154_3461_ngat) );
INVXL U_g5402 (.A(G6301_3490_gat), .Y(G6301_3490_ngat) );
INVXL U_g5403 (.A(G6308_2647_gat), .Y(G6308_2647_ngat) );
INVXL U_g5404 (.A(G5563_3481_gat), .Y(G5563_3481_ngat) );
INVXL U_g5405 (.A(G5570_2376_gat), .Y(G5570_2376_ngat) );
INVXL U_g5406 (.A(G5505_3480_gat), .Y(G5505_3480_ngat) );
INVXL U_g5407 (.A(G5512_2377_gat), .Y(G5512_2377_ngat) );
INVXL U_g5408 (.A(G5624_2076_gat), .Y(G5624_2076_ngat) );
INVXL U_g5409 (.A(G5627_3485_gat), .Y(G5627_3485_ngat) );
INVXL U_g5410 (.A(G5712_2077_gat), .Y(G5712_2077_ngat) );
INVXL U_g5411 (.A(G5715_3484_gat), .Y(G5715_3484_ngat) );
INVXL U_g5412 (.A(G5054_2121_gat), .Y(G5054_2121_ngat) );
INVXL U_g5413 (.A(G5057_3489_gat), .Y(G5057_3489_ngat) );
INVXL U_g5414 (.A(G5142_2123_gat), .Y(G5142_2123_ngat) );
INVXL U_g5415 (.A(G5145_3488_gat), .Y(G5145_3488_ngat) );
INVXL U_g5416 (.A(G6211_3491_gat), .Y(G6211_3491_ngat) );
INVXL U_g5417 (.A(G6212_3473_gat), .Y(G6212_3473_ngat) );
INVXL U_g5418 (.A(G7023_3493_gat), .Y(G7023_3493_ngat) );
INVXL U_g5419 (.A(G7030_2554_gat), .Y(G7030_2554_ngat) );
INVXL U_g5420 (.A(G6965_3492_gat), .Y(G6965_3492_ngat) );
INVXL U_g5421 (.A(G6972_2555_gat), .Y(G6972_2555_ngat) );
INVXL U_g5422 (.A(G7084_2290_gat), .Y(G7084_2290_ngat) );
INVXL U_g5423 (.A(G7087_3497_gat), .Y(G7087_3497_ngat) );
INVXL U_g5424 (.A(G7172_2291_gat), .Y(G7172_2291_ngat) );
INVXL U_g5425 (.A(G7175_3496_gat), .Y(G7175_3496_ngat) );
INVXL U_g5426 (.A(G6155_3499_gat), .Y(G6155_3499_ngat) );
INVXL U_g5427 (.A(G6162_2604_gat), .Y(G6162_2604_ngat) );
INVXL U_g5428 (.A(G6097_3498_gat), .Y(G6097_3498_ngat) );
INVXL U_g5429 (.A(G6104_2605_gat), .Y(G6104_2605_ngat) );
INVXL U_g5430 (.A(G6213_3510_gat), .Y(G6213_3510_ngat) );
INVXL U_g5431 (.A(G6220_2646_gat), .Y(G6220_2646_ngat) );
INVXL U_g5432 (.A(G6304_2370_gat), .Y(G6304_2370_ngat) );
INVXL U_g5433 (.A(G6307_3509_gat), .Y(G6307_3509_ngat) );
INVXL U_g5434 (.A(G5566_2000_gat), .Y(G5566_2000_ngat) );
INVXL U_g5435 (.A(G5569_3504_gat), .Y(G5569_3504_ngat) );
INVXL U_g5436 (.A(G5508_2001_gat), .Y(G5508_2001_ngat) );
INVXL U_g5437 (.A(G5511_3503_gat), .Y(G5511_3503_ngat) );
INVXL U_g5438 (.A(G5629_3505_gat), .Y(G5629_3505_ngat) );
INVXL U_g5439 (.A(G5630_3482_gat), .Y(G5630_3482_ngat) );
INVXL U_g5440 (.A(G5717_3506_gat), .Y(G5717_3506_ngat) );
INVXL U_g5441 (.A(G5718_3483_gat), .Y(G5718_3483_ngat) );
INVXL U_g5442 (.A(G5059_3507_gat), .Y(G5059_3507_ngat) );
INVXL U_g5443 (.A(G5060_3486_gat), .Y(G5060_3486_ngat) );
INVXL U_g5444 (.A(G5147_3508_gat), .Y(G5147_3508_ngat) );
INVXL U_g5445 (.A(G5148_3487_gat), .Y(G5148_3487_ngat) );
INVXL U_g5446 (.A(G7026_2225_gat), .Y(G7026_2225_ngat) );
INVXL U_g5447 (.A(G7029_3514_gat), .Y(G7029_3514_ngat) );
INVXL U_g5448 (.A(G6968_2226_gat), .Y(G6968_2226_ngat) );
INVXL U_g5449 (.A(G6971_3513_gat), .Y(G6971_3513_ngat) );
INVXL U_g5450 (.A(G7089_3515_gat), .Y(G7089_3515_ngat) );
INVXL U_g5451 (.A(G7090_3494_gat), .Y(G7090_3494_ngat) );
INVXL U_g5452 (.A(G7177_3516_gat), .Y(G7177_3516_ngat) );
INVXL U_g5453 (.A(G7178_3495_gat), .Y(G7178_3495_ngat) );
INVXL U_g5454 (.A(G6158_2308_gat), .Y(G6158_2308_ngat) );
INVXL U_g5455 (.A(G6161_3520_gat), .Y(G6161_3520_ngat) );
INVXL U_g5456 (.A(G6100_2309_gat), .Y(G6100_2309_ngat) );
INVXL U_g5457 (.A(G6103_3519_gat), .Y(G6103_3519_ngat) );
INVXL U_g5458 (.A(G6216_2369_gat), .Y(G6216_2369_ngat) );
INVXL U_g5459 (.A(G6219_3529_gat), .Y(G6219_3529_ngat) );
INVXL U_g5460 (.A(G6309_3522_gat), .Y(G6309_3522_ngat) );
INVXL U_g5461 (.A(G6310_3500_gat), .Y(G6310_3500_ngat) );
INVXL U_g5462 (.A(G5571_3523_gat), .Y(G5571_3523_ngat) );
INVXL U_g5463 (.A(G5572_3501_gat), .Y(G5572_3501_ngat) );
INVXL U_g5464 (.A(G5513_3524_gat), .Y(G5513_3524_ngat) );
INVXL U_g5465 (.A(G5514_3502_gat), .Y(G5514_3502_ngat) );
INVXL U_g5466 (.A(G5719_3526_gat), .Y(G5719_3526_ngat) );
INVXL U_g5467 (.A(G5726_2408_gat), .Y(G5726_2408_ngat) );
INVXL U_g5468 (.A(G5631_3525_gat), .Y(G5631_3525_ngat) );
INVXL U_g5469 (.A(G5638_2409_gat), .Y(G5638_2409_ngat) );
INVXL U_g5470 (.A(G5149_3528_gat), .Y(G5149_3528_ngat) );
INVXL U_g5471 (.A(G5156_2439_gat), .Y(G5156_2439_ngat) );
INVXL U_g5472 (.A(G5061_3527_gat), .Y(G5061_3527_ngat) );
INVXL U_g5473 (.A(G5068_2440_gat), .Y(G5068_2440_ngat) );
INVXL U_g5474 (.A(G7031_3530_gat), .Y(G7031_3530_ngat) );
INVXL U_g5475 (.A(G7032_3511_gat), .Y(G7032_3511_ngat) );
INVXL U_g5476 (.A(G6973_3531_gat), .Y(G6973_3531_ngat) );
INVXL U_g5477 (.A(G6974_3512_gat), .Y(G6974_3512_ngat) );
INVXL U_g5478 (.A(G7179_3533_gat), .Y(G7179_3533_ngat) );
INVXL U_g5479 (.A(G7186_2580_gat), .Y(G7186_2580_ngat) );
INVXL U_g5480 (.A(G7091_3532_gat), .Y(G7091_3532_ngat) );
INVXL U_g5481 (.A(G7098_2581_gat), .Y(G7098_2581_ngat) );
INVXL U_g5482 (.A(G6163_3534_gat), .Y(G6163_3534_ngat) );
INVXL U_g5483 (.A(G6164_3517_gat), .Y(G6164_3517_ngat) );
INVXL U_g5484 (.A(G6105_3535_gat), .Y(G6105_3535_ngat) );
INVXL U_g5485 (.A(G6106_3518_gat), .Y(G6106_3518_ngat) );
INVXL U_g5486 (.A(G6311_3537_gat), .Y(G6311_3537_ngat) );
INVXL U_g5487 (.A(G6318_2632_gat), .Y(G6318_2632_ngat) );
INVXL U_g5488 (.A(G6221_3536_gat), .Y(G6221_3536_ngat) );
INVXL U_g5489 (.A(G6222_3521_gat), .Y(G6222_3521_ngat) );
INVXL U_g5490 (.A(G5515_3539_gat), .Y(G5515_3539_ngat) );
INVXL U_g5491 (.A(G5522_2389_gat), .Y(G5522_2389_ngat) );
INVXL U_g5492 (.A(G5573_3538_gat), .Y(G5573_3538_ngat) );
INVXL U_g5493 (.A(G5580_2390_gat), .Y(G5580_2390_ngat) );
INVXL U_g5494 (.A(G5722_2044_gat), .Y(G5722_2044_ngat) );
INVXL U_g5495 (.A(G5725_3543_gat), .Y(G5725_3543_ngat) );
INVXL U_g5496 (.A(G5634_2045_gat), .Y(G5634_2045_ngat) );
INVXL U_g5497 (.A(G5637_3542_gat), .Y(G5637_3542_ngat) );
INVXL U_g5498 (.A(G5152_2098_gat), .Y(G5152_2098_ngat) );
INVXL U_g5499 (.A(G5155_3547_gat), .Y(G5155_3547_ngat) );
INVXL U_g5500 (.A(G5064_2099_gat), .Y(G5064_2099_ngat) );
INVXL U_g5501 (.A(G5067_3546_gat), .Y(G5067_3546_ngat) );
INVXL U_g5502 (.A(G6975_3549_gat), .Y(G6975_3549_ngat) );
INVXL U_g5503 (.A(G6982_2565_gat), .Y(G6982_2565_ngat) );
INVXL U_g5504 (.A(G7033_3548_gat), .Y(G7033_3548_ngat) );
INVXL U_g5505 (.A(G7040_2566_gat), .Y(G7040_2566_ngat) );
INVXL U_g5506 (.A(G7182_2262_gat), .Y(G7182_2262_ngat) );
INVXL U_g5507 (.A(G7185_3553_gat), .Y(G7185_3553_ngat) );
INVXL U_g5508 (.A(G7094_2263_gat), .Y(G7094_2263_ngat) );
INVXL U_g5509 (.A(G7097_3552_gat), .Y(G7097_3552_ngat) );
INVXL U_g5510 (.A(G6107_3555_gat), .Y(G6107_3555_ngat) );
INVXL U_g5511 (.A(G6114_2615_gat), .Y(G6114_2615_ngat) );
INVXL U_g5512 (.A(G6165_3554_gat), .Y(G6165_3554_ngat) );
INVXL U_g5513 (.A(G6172_2616_gat), .Y(G6172_2616_ngat) );
INVXL U_g5514 (.A(G6314_2346_gat), .Y(G6314_2346_ngat) );
INVXL U_g5515 (.A(G6317_3558_gat), .Y(G6317_3558_ngat) );
INVXL U_g5516 (.A(G6223_3557_gat), .Y(G6223_3557_ngat) );
INVXL U_g5517 (.A(G6230_2633_gat), .Y(G6230_2633_ngat) );
INVXL U_g5518 (.A(G5518_2011_gat), .Y(G5518_2011_ngat) );
INVXL U_g5519 (.A(G5521_3560_gat), .Y(G5521_3560_ngat) );
INVXL U_g5520 (.A(G5576_2013_gat), .Y(G5576_2013_ngat) );
INVXL U_g5521 (.A(G5579_3559_gat), .Y(G5579_3559_ngat) );
INVXL U_g5522 (.A(G5727_3563_gat), .Y(G5727_3563_ngat) );
INVXL U_g5523 (.A(G5728_3540_gat), .Y(G5728_3540_ngat) );
INVXL U_g5524 (.A(G5639_3564_gat), .Y(G5639_3564_ngat) );
INVXL U_g5525 (.A(G5640_3541_gat), .Y(G5640_3541_ngat) );
INVXL U_g5526 (.A(G5157_3565_gat), .Y(G5157_3565_ngat) );
INVXL U_g5527 (.A(G5158_3544_gat), .Y(G5158_3544_ngat) );
INVXL U_g5528 (.A(G5069_3566_gat), .Y(G5069_3566_ngat) );
INVXL U_g5529 (.A(G5070_3545_gat), .Y(G5070_3545_ngat) );
INVXL U_g5530 (.A(G6978_2235_gat), .Y(G6978_2235_ngat) );
INVXL U_g5531 (.A(G6981_3568_gat), .Y(G6981_3568_ngat) );
INVXL U_g5532 (.A(G7036_2237_gat), .Y(G7036_2237_ngat) );
INVXL U_g5533 (.A(G7039_3567_gat), .Y(G7039_3567_ngat) );
INVXL U_g5534 (.A(G7187_3571_gat), .Y(G7187_3571_ngat) );
INVXL U_g5535 (.A(G7188_3550_gat), .Y(G7188_3550_ngat) );
INVXL U_g5536 (.A(G7099_3572_gat), .Y(G7099_3572_ngat) );
INVXL U_g5537 (.A(G7100_3551_gat), .Y(G7100_3551_ngat) );
INVXL U_g5538 (.A(G6110_2318_gat), .Y(G6110_2318_ngat) );
INVXL U_g5539 (.A(G6113_3574_gat), .Y(G6113_3574_ngat) );
INVXL U_g5540 (.A(G6168_2320_gat), .Y(G6168_2320_ngat) );
INVXL U_g5541 (.A(G6171_3573_gat), .Y(G6171_3573_ngat) );
INVXL U_g5542 (.A(G6319_3577_gat), .Y(G6319_3577_ngat) );
INVXL U_g5543 (.A(G6320_3556_gat), .Y(G6320_3556_ngat) );
INVXL U_g5544 (.A(G6226_2347_gat), .Y(G6226_2347_ngat) );
INVXL U_g5545 (.A(G6229_3579_gat), .Y(G6229_3579_ngat) );
INVXL U_g5546 (.A(G1755_3580_gat), .Y(G1755_3580_ngat) );
INVXL U_g5547 (.A(G1756_3561_gat), .Y(G1756_3561_ngat) );
INVXL U_g5548 (.A(G1760_3581_gat), .Y(G1760_3581_ngat) );
INVXL U_g5549 (.A(G1761_3562_gat), .Y(G1761_3562_ngat) );
INVXL U_g5550 (.A(G5729_3582_gat), .Y(G5729_3582_ngat) );
INVXL U_g5551 (.A(G5736_2421_gat), .Y(G5736_2421_ngat) );
INVXL U_g5552 (.A(G5641_3583_gat), .Y(G5641_3583_ngat) );
INVXL U_g5553 (.A(G5648_2422_gat), .Y(G5648_2422_ngat) );
INVXL U_g5554 (.A(G5159_3584_gat), .Y(G5159_3584_ngat) );
INVXL U_g5555 (.A(G5166_2483_gat), .Y(G5166_2483_ngat) );
INVXL U_g5556 (.A(G5071_3585_gat), .Y(G5071_3585_ngat) );
INVXL U_g5557 (.A(G5078_2484_gat), .Y(G5078_2484_ngat) );
INVXL U_g5558 (.A(G4057_3586_gat), .Y(G4057_3586_ngat) );
INVXL U_g5559 (.A(G4058_3569_gat), .Y(G4058_3569_ngat) );
INVXL U_g5560 (.A(G4062_3587_gat), .Y(G4062_3587_ngat) );
INVXL U_g5561 (.A(G4063_3570_gat), .Y(G4063_3570_ngat) );
INVXL U_g5562 (.A(G7189_3588_gat), .Y(G7189_3588_ngat) );
INVXL U_g5563 (.A(G7196_2591_gat), .Y(G7196_2591_ngat) );
INVXL U_g5564 (.A(G7101_3589_gat), .Y(G7101_3589_ngat) );
INVXL U_g5565 (.A(G7108_2592_gat), .Y(G7108_2592_ngat) );
INVXL U_g5566 (.A(G2817_3590_gat), .Y(G2817_3590_ngat) );
INVXL U_g5567 (.A(G2818_3575_gat), .Y(G2818_3575_ngat) );
INVXL U_g5568 (.A(G2822_3591_gat), .Y(G2822_3591_ngat) );
INVXL U_g5569 (.A(G2823_3576_gat), .Y(G2823_3576_ngat) );
INVXL U_g5570 (.A(G6231_3593_gat), .Y(G6231_3593_ngat) );
INVXL U_g5571 (.A(G6232_3578_gat), .Y(G6232_3578_ngat) );
INVXL U_g5572 (.A(G6321_3592_gat), .Y(G6321_3592_ngat) );
INVXL U_g5573 (.A(G6328_2642_gat), .Y(G6328_2642_ngat) );
INVXL U_g5574 (.A(G5732_2063_gat), .Y(G5732_2063_ngat) );
INVXL U_g5575 (.A(G5735_3596_gat), .Y(G5735_3596_ngat) );
INVXL U_g5576 (.A(G5644_2064_gat), .Y(G5644_2064_ngat) );
INVXL U_g5577 (.A(G5647_3597_gat), .Y(G5647_3597_ngat) );
INVXL U_g5578 (.A(G5162_2166_gat), .Y(G5162_2166_ngat) );
INVXL U_g5579 (.A(G5165_3600_gat), .Y(G5165_3600_ngat) );
INVXL U_g5580 (.A(G5074_2167_gat), .Y(G5074_2167_ngat) );
INVXL U_g5581 (.A(G5077_3601_gat), .Y(G5077_3601_ngat) );
INVXL U_g5582 (.A(G7192_2278_gat), .Y(G7192_2278_ngat) );
INVXL U_g5583 (.A(G7195_3606_gat), .Y(G7195_3606_ngat) );
INVXL U_g5584 (.A(G7104_2279_gat), .Y(G7104_2279_ngat) );
INVXL U_g5585 (.A(G7107_3607_gat), .Y(G7107_3607_ngat) );
INVXL U_g5586 (.A(G6324_2359_gat), .Y(G6324_2359_ngat) );
INVXL U_g5587 (.A(G6327_3612_gat), .Y(G6327_3612_ngat) );
INVXL U_g5588 (.A(G6233_3613_gat), .Y(G6233_3613_ngat) );
INVXL U_g5589 (.A(G6240_2643_gat), .Y(G6240_2643_ngat) );
INVXL U_g5590 (.A(G5659_3619_gat), .Y(G5659_3619_ngat) );
INVXL U_g5591 (.A(G5660_3598_gat), .Y(G5660_3598_ngat) );
INVXL U_g5592 (.A(G5649_3620_gat), .Y(G5649_3620_ngat) );
INVXL U_g5593 (.A(G5650_3599_gat), .Y(G5650_3599_ngat) );
INVXL U_g5594 (.A(G5089_3621_gat), .Y(G5089_3621_ngat) );
INVXL U_g5595 (.A(G5090_3602_gat), .Y(G5090_3602_ngat) );
INVXL U_g5596 (.A(G5079_3622_gat), .Y(G5079_3622_ngat) );
INVXL U_g5597 (.A(G5080_3603_gat), .Y(G5080_3603_ngat) );
INVXL U_g5598 (.A(G7119_3631_gat), .Y(G7119_3631_ngat) );
INVXL U_g5599 (.A(G7120_3608_gat), .Y(G7120_3608_ngat) );
INVXL U_g5600 (.A(G7109_3632_gat), .Y(G7109_3632_ngat) );
INVXL U_g5601 (.A(G7110_3609_gat), .Y(G7110_3609_ngat) );
INVXL U_g5602 (.A(G6251_3634_gat), .Y(G6251_3634_ngat) );
INVXL U_g5603 (.A(G6252_3614_gat), .Y(G6252_3614_ngat) );
INVXL U_g5604 (.A(G6236_2360_gat), .Y(G6236_2360_ngat) );
INVXL U_g5605 (.A(G6239_3633_gat), .Y(G6239_3633_ngat) );
INVXL U_g5606 (.A(G5661_3637_gat), .Y(G5661_3637_ngat) );
INVXL U_g5607 (.A(G5668_2416_gat), .Y(G5668_2416_ngat) );
INVXL U_g5608 (.A(G5651_3638_gat), .Y(G5651_3638_ngat) );
INVXL U_g5609 (.A(G5658_2417_gat), .Y(G5658_2417_ngat) );
INVXL U_g5610 (.A(G5091_3639_gat), .Y(G5091_3639_ngat) );
INVXL U_g5611 (.A(G5098_2446_gat), .Y(G5098_2446_ngat) );
INVXL U_g5612 (.A(G5081_3640_gat), .Y(G5081_3640_ngat) );
INVXL U_g5613 (.A(G5088_2447_gat), .Y(G5088_2447_ngat) );
INVXL U_g5614 (.A(G7121_3643_gat), .Y(G7121_3643_ngat) );
INVXL U_g5615 (.A(G7128_2587_gat), .Y(G7128_2587_ngat) );
INVXL U_g5616 (.A(G7111_3644_gat), .Y(G7111_3644_ngat) );
INVXL U_g5617 (.A(G7118_2588_gat), .Y(G7118_2588_ngat) );
INVXL U_g5618 (.A(G6253_3645_gat), .Y(G6253_3645_ngat) );
INVXL U_g5619 (.A(G6260_2636_gat), .Y(G6260_2636_ngat) );
INVXL U_g5620 (.A(G6241_3646_gat), .Y(G6241_3646_ngat) );
INVXL U_g5621 (.A(G6242_3635_gat), .Y(G6242_3635_ngat) );
INVXL U_g5622 (.A(G5664_2052_gat), .Y(G5664_2052_ngat) );
INVXL U_g5623 (.A(G5667_3650_gat), .Y(G5667_3650_ngat) );
INVXL U_g5624 (.A(G5654_2054_gat), .Y(G5654_2054_ngat) );
INVXL U_g5625 (.A(G5657_3651_gat), .Y(G5657_3651_ngat) );
INVXL U_g5626 (.A(G5094_2106_gat), .Y(G5094_2106_ngat) );
INVXL U_g5627 (.A(G5097_3654_gat), .Y(G5097_3654_ngat) );
INVXL U_g5628 (.A(G5084_2108_gat), .Y(G5084_2108_ngat) );
INVXL U_g5629 (.A(G5087_3655_gat), .Y(G5087_3655_ngat) );
INVXL U_g5630 (.A(G7124_2270_gat), .Y(G7124_2270_ngat) );
INVXL U_g5631 (.A(G7127_3660_gat), .Y(G7127_3660_ngat) );
INVXL U_g5632 (.A(G7114_2272_gat), .Y(G7114_2272_ngat) );
INVXL U_g5633 (.A(G7117_3661_gat), .Y(G7117_3661_ngat) );
INVXL U_g5634 (.A(G6256_2350_gat), .Y(G6256_2350_ngat) );
INVXL U_g5635 (.A(G6259_3663_gat), .Y(G6259_3663_ngat) );
INVXL U_g5636 (.A(G6243_3664_gat), .Y(G6243_3664_ngat) );
INVXL U_g5637 (.A(G6250_2638_gat), .Y(G6250_2638_ngat) );
INVXL U_g5638 (.A(G1778_3665_gat), .Y(G1778_3665_ngat) );
INVXL U_g5639 (.A(G1779_3648_gat), .Y(G1779_3648_ngat) );
INVXL U_g5640 (.A(G1775_3666_gat), .Y(G1775_3666_ngat) );
INVXL U_g5641 (.A(G1776_3649_gat), .Y(G1776_3649_ngat) );
INVXL U_g5642 (.A(G987_3667_gat), .Y(G987_3667_ngat) );
INVXL U_g5643 (.A(G988_3652_gat), .Y(G988_3652_ngat) );
INVXL U_g5644 (.A(G984_3668_gat), .Y(G984_3668_ngat) );
INVXL U_g5645 (.A(G985_3653_gat), .Y(G985_3653_ngat) );
INVXL U_g5646 (.A(G4079_3669_gat), .Y(G4079_3669_ngat) );
INVXL U_g5647 (.A(G4080_3658_gat), .Y(G4080_3658_ngat) );
INVXL U_g5648 (.A(G4076_3670_gat), .Y(G4076_3670_ngat) );
INVXL U_g5649 (.A(G4077_3659_gat), .Y(G4077_3659_ngat) );
INVXL U_g5650 (.A(G2840_3671_gat), .Y(G2840_3671_ngat) );
INVXL U_g5651 (.A(G2841_3662_gat), .Y(G2841_3662_ngat) );
INVXL U_g5652 (.A(G6246_2351_gat), .Y(G6246_2351_ngat) );
INVXL U_g5653 (.A(G6249_3673_gat), .Y(G6249_3673_ngat) );
INVXL U_g5654 (.A(G2837_3682_gat), .Y(G2837_3682_ngat) );
INVXL U_g5655 (.A(G2838_3672_gat), .Y(G2838_3672_ngat) );
INVXL U_g5656 (.A(G5740_3694_gat), .Y(G5740_3694_ngat) );
INVXL U_g5657 (.A(G5743_3647_gat), .Y(G5743_3647_ngat) );
INVXL U_g5658 (.A(G5170_3696_gat), .Y(G5170_3696_ngat) );
INVXL U_g5659 (.A(G5173_3469_gat), .Y(G5173_3469_ngat) );
INVXL U_g5660 (.A(G6332_3697_gat), .Y(G6332_3697_ngat) );
INVXL U_g5661 (.A(G6335_3656_gat), .Y(G6335_3656_ngat) );
INVXL U_g5662 (.A(G7200_3699_gat), .Y(G7200_3699_ngat) );
INVXL U_g5663 (.A(G7203_3657_gat), .Y(G7203_3657_ngat) );
INVXL U_g5664 (.A(G5737_3636_gat), .Y(G5737_3636_ngat) );
INVXL U_g5665 (.A(G5744_3698_gat), .Y(G5744_3698_ngat) );
INVXL U_g5666 (.A(G5167_3446_gat), .Y(G5167_3446_ngat) );
INVXL U_g5667 (.A(G5174_3700_gat), .Y(G5174_3700_ngat) );
INVXL U_g5668 (.A(G6329_3641_gat), .Y(G6329_3641_ngat) );
INVXL U_g5669 (.A(G6336_3704_gat), .Y(G6336_3704_ngat) );
INVXL U_g5670 (.A(G7197_3642_gat), .Y(G7197_3642_ngat) );
INVXL U_g5671 (.A(G7204_3706_gat), .Y(G7204_3706_ngat) );
INVXL U_g5672 (.A(G1791_3701_gat), .Y(G1791_3701_ngat) );
INVXL U_g5673 (.A(G1792_3707_gat), .Y(G1792_3707_ngat) );
INVXL U_g5674 (.A(G1003_3702_gat), .Y(G1003_3702_ngat) );
INVXL U_g5675 (.A(G1004_3708_gat), .Y(G1004_3708_ngat) );
INVXL U_g5676 (.A(G2855_3703_gat), .Y(G2855_3703_ngat) );
INVXL U_g5677 (.A(G2856_3709_gat), .Y(G2856_3709_ngat) );
INVXL U_g5678 (.A(G4092_3705_gat), .Y(G4092_3705_ngat) );
INVXL U_g5679 (.A(G4093_3710_gat), .Y(G4093_3710_ngat) );

endmodule
