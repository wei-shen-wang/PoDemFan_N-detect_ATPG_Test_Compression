module C5315 ( G1P0gat, G4P1gat, G11P2gat, G14P3gat, G17P4gat, G20P5gat, G23P6gat, G24P7gat, G25P8gat, G26P9gat, G27P10gat, G31P11gat, G34P12gat, G37P13gat, G40P14gat, G43P15gat, G46P16gat, G49P17gat, G52P18gat, G53P19gat, G54P20gat, G61P21gat, G64P22gat, G67P23gat, G70P24gat, G73P25gat, G76P26gat, G79P27gat, G80P28gat, G81P29gat, G82P30gat, G83P31gat, G86P32gat, G87P33gat, G88P34gat, G91P35gat, G94P36gat, G97P37gat, G100P38gat, G103P39gat, G106P40gat, G109P41gat, G112P42gat, G113P43gat, G114P44gat, G115P45gat, G116P46gat, G117P47gat, G118P48gat, G119P49gat, G120P50gat, G121P51gat, G122P52gat, G123P53gat, G126P54gat, G127P55gat, G128P56gat, G129P57gat, G130P58gat, G131P59gat, G132P60gat, G135P61gat, G136P62gat, G137P63gat, G140P64gat, G141P65gat, G145P66gat, G146P67gat, G149P68gat, G152P69gat, G155P70gat, G158P71gat, G161P72gat, G164P73gat, G167P74gat, G170P75gat, G173P76gat, G176P77gat, G179P78gat, G182P79gat, G185P80gat, G188P81gat, G191P82gat, G194P83gat, G197P84gat, G200P85gat, G203P86gat, G206P87gat, G209P88gat, G210P89gat, G217P90gat, G218P91gat, G225P92gat, G226P93gat, G233P94gat, G234P95gat, G241P96gat, G242P97gat, G245P98gat, G248P99gat, G251P100gat, G254P101gat, G257P102gat, G264P103gat, G265P104gat, G272P105gat, G273P106gat, G280P107gat, G281P108gat, G288P109gat, G289P110gat, G292P111gat, G293P112gat, G299P113gat, G302P114gat, G307P115gat, G308P116gat, G315P117gat, G316P118gat, G323P119gat, G324P120gat, G331P121gat, G332P122gat, G335P123gat, G338P124gat, G341P125gat, G348P126gat, G351P127gat, G358P128gat, G361P129gat, G366P130gat, G369P131gat, G372P132gat, G373P133gat, G374P134gat, G386P135gat, G389P136gat, G400P137gat, G411P138gat, G422P139gat, G435P140gat, G446P141gat, G457P142gat, G468P143gat, G479P144gat, G490P145gat, G503P146gat, G514P147gat, G523P148gat, G534P149gat, G545P150gat, G549P151gat, G552P152gat, G556P153gat, G559P154gat, G562P155gat, G1497P156gat, G1689P157gat, G1690P158gat, G1691P159gat, G1694P160gat, G2174P161gat, G2358P162gat, G2824P163gat, G3173P164gat, G3546P165gat, G3548P166gat, G3550P167gat, G3552P168gat, G3717P169gat, G3724P170gat, G4087P171gat, G4088P172gat, G4089P173gat, G4090P174gat, G4091P175gat, G4092P176gat, G4115P177gat, G144P354gat, G298P299gat, G973P202gat, G594P224gat, G599P269gat, G600P259gat, G601P220gat, G602P222gat, G603P225gat, G604P223gat, G611P275gat, G612P263gat, G810P356gat, G848P330gat, G849P219gat, G850P217gat, G851P218gat, G634P665gat, G815P627gat, G845P845gat, G847P465gat, G926P624gat, G923P619gat, G921P664gat, G892P408gat, G887P528gat, G606P407gat, G656P621gat, G809P655gat, G993P850gat, G978P851gat, G949P852gat, G939P853gat, G889P734gat, G593P733gat, G636P1280gat, G704P1281gat, G717P1282gat, G820P1283gat, G639P1275gat, G673P1276gat, G707P1277gat, G715P1278gat, G598P1623gat, G610P1519gat, G588P1696gat, G615P1750gat, G626P1752gat, G632P1692gat, G1002P1920gat, G1004P1977gat, G591P1894gat, G618P1925gat, G621P1893gat, G629P1926gat, G822P1933gat, G838P2064gat, G861P2070gat, G623P2152gat, G722P2131gat, G832P2133gat, G834P2123gat, G836P2128gat, G859P2132gat, G871P2127gat, G873P2124gat, G875P2125gat, G877P2126gat, G998P2163gat, G1000P2168gat, G575P2240gat, G585P2236gat, G661P2178gat, G693P2179gat, G747P2187gat, G752P2189gat, G757P2190gat, G762P2184gat, G787P2186gat, G792P2188gat, G797P2191gat, G802P2183gat, G642P2222gat, G664P2223gat, G667P2224gat, G670P2225gat, G676P2229gat, G696P2226gat, G699P2227gat, G702P2228gat, G818P2273gat, G813P2260gat, G824P2274gat, G826P2275gat, G828P2233gat, G830P2182gat, G854P2268gat, G863P2276gat, G865P2277gat, G867P2237gat, G869P2181gat, G712P2297gat, G727P2298gat, G732P2300gat, G737P2279gat, G742P2238gat, G772P2299gat, G777P2278gat, G782P2239gat, G645P2271gat, G648P2295gat, G651P2314gat, G654P2315gat, G679P2272gat, G682P2296gat, G685P2316gat, G688P2317gat, G843P2455gat, G882P2456gat, G767P2479gat, G807P2480gat, G658P2483gat, G690P2484gat);

input G1P0gat;
input G4P1gat;
input G11P2gat;
input G14P3gat;
input G17P4gat;
input G20P5gat;
input G23P6gat;
input G24P7gat;
input G25P8gat;
input G26P9gat;
input G27P10gat;
input G31P11gat;
input G34P12gat;
input G37P13gat;
input G40P14gat;
input G43P15gat;
input G46P16gat;
input G49P17gat;
input G52P18gat;
input G53P19gat;
input G54P20gat;
input G61P21gat;
input G64P22gat;
input G67P23gat;
input G70P24gat;
input G73P25gat;
input G76P26gat;
input G79P27gat;
input G80P28gat;
input G81P29gat;
input G82P30gat;
input G83P31gat;
input G86P32gat;
input G87P33gat;
input G88P34gat;
input G91P35gat;
input G94P36gat;
input G97P37gat;
input G100P38gat;
input G103P39gat;
input G106P40gat;
input G109P41gat;
input G112P42gat;
input G113P43gat;
input G114P44gat;
input G115P45gat;
input G116P46gat;
input G117P47gat;
input G118P48gat;
input G119P49gat;
input G120P50gat;
input G121P51gat;
input G122P52gat;
input G123P53gat;
input G126P54gat;
input G127P55gat;
input G128P56gat;
input G129P57gat;
input G130P58gat;
input G131P59gat;
input G132P60gat;
input G135P61gat;
input G136P62gat;
input G137P63gat;
input G140P64gat;
input G141P65gat;
input G145P66gat;
input G146P67gat;
input G149P68gat;
input G152P69gat;
input G155P70gat;
input G158P71gat;
input G161P72gat;
input G164P73gat;
input G167P74gat;
input G170P75gat;
input G173P76gat;
input G176P77gat;
input G179P78gat;
input G182P79gat;
input G185P80gat;
input G188P81gat;
input G191P82gat;
input G194P83gat;
input G197P84gat;
input G200P85gat;
input G203P86gat;
input G206P87gat;
input G209P88gat;
input G210P89gat;
input G217P90gat;
input G218P91gat;
input G225P92gat;
input G226P93gat;
input G233P94gat;
input G234P95gat;
input G241P96gat;
input G242P97gat;
input G245P98gat;
input G248P99gat;
input G251P100gat;
input G254P101gat;
input G257P102gat;
input G264P103gat;
input G265P104gat;
input G272P105gat;
input G273P106gat;
input G280P107gat;
input G281P108gat;
input G288P109gat;
input G289P110gat;
input G292P111gat;
input G293P112gat;
input G299P113gat;
input G302P114gat;
input G307P115gat;
input G308P116gat;
input G315P117gat;
input G316P118gat;
input G323P119gat;
input G324P120gat;
input G331P121gat;
input G332P122gat;
input G335P123gat;
input G338P124gat;
input G341P125gat;
input G348P126gat;
input G351P127gat;
input G358P128gat;
input G361P129gat;
input G366P130gat;
input G369P131gat;
input G372P132gat;
input G373P133gat;
input G374P134gat;
input G386P135gat;
input G389P136gat;
input G400P137gat;
input G411P138gat;
input G422P139gat;
input G435P140gat;
input G446P141gat;
input G457P142gat;
input G468P143gat;
input G479P144gat;
input G490P145gat;
input G503P146gat;
input G514P147gat;
input G523P148gat;
input G534P149gat;
input G545P150gat;
input G549P151gat;
input G552P152gat;
input G556P153gat;
input G559P154gat;
input G562P155gat;
input G1497P156gat;
input G1689P157gat;
input G1690P158gat;
input G1691P159gat;
input G1694P160gat;
input G2174P161gat;
input G2358P162gat;
input G2824P163gat;
input G3173P164gat;
input G3546P165gat;
input G3548P166gat;
input G3550P167gat;
input G3552P168gat;
input G3717P169gat;
input G3724P170gat;
input G4087P171gat;
input G4088P172gat;
input G4089P173gat;
input G4090P174gat;
input G4091P175gat;
input G4092P176gat;
input G4115P177gat;

output G144P354gat;
output G298P299gat;
output G973P202gat;
output G594P224gat;
output G599P269gat;
output G600P259gat;
output G601P220gat;
output G602P222gat;
output G603P225gat;
output G604P223gat;
output G611P275gat;
output G612P263gat;
output G810P356gat;
output G848P330gat;
output G849P219gat;
output G850P217gat;
output G851P218gat;
output G634P665gat;
output G815P627gat;
output G845P845gat;
output G847P465gat;
output G926P624gat;
output G923P619gat;
output G921P664gat;
output G892P408gat;
output G887P528gat;
output G606P407gat;
output G656P621gat;
output G809P655gat;
output G993P850gat;
output G978P851gat;
output G949P852gat;
output G939P853gat;
output G889P734gat;
output G593P733gat;
output G636P1280gat;
output G704P1281gat;
output G717P1282gat;
output G820P1283gat;
output G639P1275gat;
output G673P1276gat;
output G707P1277gat;
output G715P1278gat;
output G598P1623gat;
output G610P1519gat;
output G588P1696gat;
output G615P1750gat;
output G626P1752gat;
output G632P1692gat;
output G1002P1920gat;
output G1004P1977gat;
output G591P1894gat;
output G618P1925gat;
output G621P1893gat;
output G629P1926gat;
output G822P1933gat;
output G838P2064gat;
output G861P2070gat;
output G623P2152gat;
output G722P2131gat;
output G832P2133gat;
output G834P2123gat;
output G836P2128gat;
output G859P2132gat;
output G871P2127gat;
output G873P2124gat;
output G875P2125gat;
output G877P2126gat;
output G998P2163gat;
output G1000P2168gat;
output G575P2240gat;
output G585P2236gat;
output G661P2178gat;
output G693P2179gat;
output G747P2187gat;
output G752P2189gat;
output G757P2190gat;
output G762P2184gat;
output G787P2186gat;
output G792P2188gat;
output G797P2191gat;
output G802P2183gat;
output G642P2222gat;
output G664P2223gat;
output G667P2224gat;
output G670P2225gat;
output G676P2229gat;
output G696P2226gat;
output G699P2227gat;
output G702P2228gat;
output G818P2273gat;
output G813P2260gat;
output G824P2274gat;
output G826P2275gat;
output G828P2233gat;
output G830P2182gat;
output G854P2268gat;
output G863P2276gat;
output G865P2277gat;
output G867P2237gat;
output G869P2181gat;
output G712P2297gat;
output G727P2298gat;
output G732P2300gat;
output G737P2279gat;
output G742P2238gat;
output G772P2299gat;
output G777P2278gat;
output G782P2239gat;
output G645P2271gat;
output G648P2295gat;
output G651P2314gat;
output G654P2315gat;
output G679P2272gat;
output G682P2296gat;
output G685P2316gat;
output G688P2317gat;
output G843P2455gat;
output G882P2456gat;
output G767P2479gat;
output G807P2480gat;
output G658P2483gat;
output G690P2484gat;

BUFX20 U_g144P354 (.A(G141P65gat), .Y(G144P354gat) );
BUFX20 U_g298P299 (.A(G293P112gat), .Y(G298P299gat) );
BUFX20 U_g973P202 (.A(G3173P164gat), .Y(G973P202gat) );
BUFX20 U_g594P224 (.A(GB3gat), .Y(G594P224gat) );
BUFX20 U_g599P269 (.A(GB4gat), .Y(G599P269gat) );
BUFX20 U_g600P259 (.A(GB5gat), .Y(G600P259gat) );
BUFX20 U_g601P220 (.A(GB6gat), .Y(G601P220gat) );
BUFX20 U_g602P222 (.A(GB7gat), .Y(G602P222gat) );
BUFX20 U_g603P225 (.A(GB8gat), .Y(G603P225gat) );
BUFX20 U_g604P223 (.A(GB9gat), .Y(G604P223gat) );
BUFX20 U_g611P275 (.A(GB10gat), .Y(G611P275gat) );
BUFX20 U_g612P263 (.A(GB11gat), .Y(G612P263gat) );
BUFX20 U_g810P356 (.A(GB12gat), .Y(G810P356gat) );
BUFX20 U_g848P330 (.A(GB13gat), .Y(G848P330gat) );
BUFX20 U_g849P219 (.A(GB14gat), .Y(G849P219gat) );
BUFX20 U_g850P217 (.A(GB15gat), .Y(G850P217gat) );
BUFX20 U_g851P218 (.A(GB16gat), .Y(G851P218gat) );
BUFX20 U_g634P665 (.A(GB17gat), .Y(G634P665gat) );
BUFX20 U_g815P627 (.A(GB18gat), .Y(G815P627gat) );
BUFX20 U_g845P845 (.A(GB19gat), .Y(G845P845gat) );
BUFX20 U_g847P465 (.A(GB20gat), .Y(G847P465gat) );
BUFX20 U_g926P624 (.A(G137P63gat), .Y(G926P624gat) );
BUFX20 U_g923P619 (.A(G141P65gat), .Y(G923P619gat) );
BUFX20 U_g921P664 (.A(G1P0gat), .Y(G921P664gat) );
BUFX20 U_g892P408 (.A(G549P151gat), .Y(G892P408gat) );
BUFX20 U_g887P528 (.A(G299P113gat), .Y(G887P528gat) );
BUFX20 U_g606P407 (.A(GB26gat), .Y(G606P407gat) );
BUFX20 U_g656P621 (.A(GB27gat), .Y(G656P621gat) );
BUFX20 U_g809P655 (.A(GB28gat), .Y(G809P655gat) );
BUFX20 U_g993P850 (.A(G1P0gat), .Y(G993P850gat) );
BUFX20 U_g978P851 (.A(G1P0gat), .Y(G978P851gat) );
BUFX20 U_g949P852 (.A(G1P0gat), .Y(G949P852gat) );
BUFX20 U_g939P853 (.A(G1P0gat), .Y(G939P853gat) );
BUFX20 U_g889P734 (.A(G299P113gat), .Y(G889P734gat) );
BUFX20 U_g593P733 (.A(GB34gat), .Y(G593P733gat) );
BUFX20 U_g636P1280 (.A(GB35gat), .Y(G636P1280gat) );
BUFX20 U_g704P1281 (.A(GB36gat), .Y(G704P1281gat) );
BUFX20 U_g717P1282 (.A(GB37gat), .Y(G717P1282gat) );
BUFX20 U_g820P1283 (.A(GB38gat), .Y(G820P1283gat) );
BUFX20 U_g639P1275 (.A(GB39gat), .Y(G639P1275gat) );
BUFX20 U_g673P1276 (.A(GB40gat), .Y(G673P1276gat) );
BUFX20 U_g707P1277 (.A(GB41gat), .Y(G707P1277gat) );
BUFX20 U_g715P1278 (.A(GB42gat), .Y(G715P1278gat) );
BUFX20 U_g598P1623 (.A(GB43gat), .Y(G598P1623gat) );
BUFX20 U_g610P1519 (.A(GB44gat), .Y(G610P1519gat) );
BUFX20 U_g588P1696 (.A(GB45gat), .Y(G588P1696gat) );
BUFX20 U_g615P1750 (.A(GB46gat), .Y(G615P1750gat) );
BUFX20 U_g626P1752 (.A(GB47gat), .Y(G626P1752gat) );
BUFX20 U_g632P1692 (.A(GB48gat), .Y(G632P1692gat) );
BUFX20 U_g1002P1920 (.A(GB49gat), .Y(G1002P1920gat) );
BUFX20 U_g1004P1977 (.A(GB50gat), .Y(G1004P1977gat) );
BUFX20 U_g591P1894 (.A(GB51gat), .Y(G591P1894gat) );
BUFX20 U_g618P1925 (.A(GB52gat), .Y(G618P1925gat) );
BUFX20 U_g621P1893 (.A(GB53gat), .Y(G621P1893gat) );
BUFX20 U_g629P1926 (.A(GB54gat), .Y(G629P1926gat) );
BUFX20 U_g822P1933 (.A(GB55gat), .Y(G822P1933gat) );
BUFX20 U_g838P2064 (.A(GB56gat), .Y(G838P2064gat) );
BUFX20 U_g861P2070 (.A(GB57gat), .Y(G861P2070gat) );
BUFX20 U_g623P2152 (.A(GB58gat), .Y(G623P2152gat) );
BUFX20 U_g722P2131 (.A(GB59gat), .Y(G722P2131gat) );
BUFX20 U_g832P2133 (.A(GB60gat), .Y(G832P2133gat) );
BUFX20 U_g834P2123 (.A(GB61gat), .Y(G834P2123gat) );
BUFX20 U_g836P2128 (.A(GB62gat), .Y(G836P2128gat) );
BUFX20 U_g859P2132 (.A(GB63gat), .Y(G859P2132gat) );
BUFX20 U_g871P2127 (.A(GB64gat), .Y(G871P2127gat) );
BUFX20 U_g873P2124 (.A(GB65gat), .Y(G873P2124gat) );
BUFX20 U_g875P2125 (.A(GB66gat), .Y(G875P2125gat) );
BUFX20 U_g877P2126 (.A(GB67gat), .Y(G877P2126gat) );
BUFX20 U_g998P2163 (.A(GB68gat), .Y(G998P2163gat) );
BUFX20 U_g1000P2168 (.A(GB69gat), .Y(G1000P2168gat) );
BUFX20 U_g575P2240 (.A(GB70gat), .Y(G575P2240gat) );
BUFX20 U_g585P2236 (.A(GB71gat), .Y(G585P2236gat) );
BUFX20 U_g661P2178 (.A(GB72gat), .Y(G661P2178gat) );
BUFX20 U_g693P2179 (.A(GB73gat), .Y(G693P2179gat) );
BUFX20 U_g747P2187 (.A(GB74gat), .Y(G747P2187gat) );
BUFX20 U_g752P2189 (.A(GB75gat), .Y(G752P2189gat) );
BUFX20 U_g757P2190 (.A(GB76gat), .Y(G757P2190gat) );
BUFX20 U_g762P2184 (.A(GB77gat), .Y(G762P2184gat) );
BUFX20 U_g787P2186 (.A(GB78gat), .Y(G787P2186gat) );
BUFX20 U_g792P2188 (.A(GB79gat), .Y(G792P2188gat) );
BUFX20 U_g797P2191 (.A(GB80gat), .Y(G797P2191gat) );
BUFX20 U_g802P2183 (.A(GB81gat), .Y(G802P2183gat) );
BUFX20 U_g642P2222 (.A(GB82gat), .Y(G642P2222gat) );
BUFX20 U_g664P2223 (.A(GB83gat), .Y(G664P2223gat) );
BUFX20 U_g667P2224 (.A(GB84gat), .Y(G667P2224gat) );
BUFX20 U_g670P2225 (.A(GB85gat), .Y(G670P2225gat) );
BUFX20 U_g676P2229 (.A(GB86gat), .Y(G676P2229gat) );
BUFX20 U_g696P2226 (.A(GB87gat), .Y(G696P2226gat) );
BUFX20 U_g699P2227 (.A(GB88gat), .Y(G699P2227gat) );
BUFX20 U_g702P2228 (.A(GB89gat), .Y(G702P2228gat) );
BUFX20 U_g818P2273 (.A(GB90gat), .Y(G818P2273gat) );
BUFX20 U_g813P2260 (.A(GB91gat), .Y(G813P2260gat) );
BUFX20 U_g824P2274 (.A(GB92gat), .Y(G824P2274gat) );
BUFX20 U_g826P2275 (.A(GB93gat), .Y(G826P2275gat) );
BUFX20 U_g828P2233 (.A(GB94gat), .Y(G828P2233gat) );
BUFX20 U_g830P2182 (.A(GB95gat), .Y(G830P2182gat) );
BUFX20 U_g854P2268 (.A(GB96gat), .Y(G854P2268gat) );
BUFX20 U_g863P2276 (.A(GB97gat), .Y(G863P2276gat) );
BUFX20 U_g865P2277 (.A(GB98gat), .Y(G865P2277gat) );
BUFX20 U_g867P2237 (.A(GB99gat), .Y(G867P2237gat) );
BUFX20 U_g869P2181 (.A(GB100gat), .Y(G869P2181gat) );
BUFX20 U_g712P2297 (.A(GB101gat), .Y(G712P2297gat) );
BUFX20 U_g727P2298 (.A(GB102gat), .Y(G727P2298gat) );
BUFX20 U_g732P2300 (.A(GB103gat), .Y(G732P2300gat) );
BUFX20 U_g737P2279 (.A(GB104gat), .Y(G737P2279gat) );
BUFX20 U_g742P2238 (.A(GB105gat), .Y(G742P2238gat) );
BUFX20 U_g772P2299 (.A(GB106gat), .Y(G772P2299gat) );
BUFX20 U_g777P2278 (.A(GB107gat), .Y(G777P2278gat) );
BUFX20 U_g782P2239 (.A(GB108gat), .Y(G782P2239gat) );
BUFX20 U_g645P2271 (.A(GB109gat), .Y(G645P2271gat) );
BUFX20 U_g648P2295 (.A(GB110gat), .Y(G648P2295gat) );
BUFX20 U_g651P2314 (.A(GB111gat), .Y(G651P2314gat) );
BUFX20 U_g654P2315 (.A(GB112gat), .Y(G654P2315gat) );
BUFX20 U_g679P2272 (.A(GB113gat), .Y(G679P2272gat) );
BUFX20 U_g682P2296 (.A(GB114gat), .Y(G682P2296gat) );
BUFX20 U_g685P2316 (.A(GB115gat), .Y(G685P2316gat) );
BUFX20 U_g688P2317 (.A(GB116gat), .Y(G688P2317gat) );
BUFX20 U_g843P2455 (.A(GB117gat), .Y(G843P2455gat) );
BUFX20 U_g882P2456 (.A(GB118gat), .Y(G882P2456gat) );
BUFX20 U_g767P2479 (.A(GB119gat), .Y(G767P2479gat) );
BUFX20 U_g807P2480 (.A(GB120gat), .Y(G807P2480gat) );
BUFX20 U_g658P2483 (.A(GB121gat), .Y(G658P2483gat) );
BUFX20 U_g690P2484 (.A(GB122gat), .Y(G690P2484gat) );
INVXL U_gB3 (.A(G545P150gat), .Y(GB3gat) );
INVXL U_gB4 (.A(G348P126gat), .Y(GB4gat) );
INVXL U_gB5 (.A(G366P130gat), .Y(GB5gat) );
AND2XL U_gB6 (.A(G552P152gat), .B(G562P155gat), .Y(GB6gat) );
INVXL U_gB7 (.A(G549P151gat), .Y(GB7gat) );
INVXL U_gB8 (.A(G545P150gat), .Y(GB8gat) );
INVXL U_gB9 (.A(G545P150gat), .Y(GB9gat) );
INVXL U_gB10 (.A(G338P124gat), .Y(GB10gat) );
INVXL U_gB11 (.A(G358P128gat), .Y(GB11gat) );
AND2XL U_gB12 (.A(G141P65gat), .B(G145P66gat), .Y(GB12gat) );
INVXL U_gB13 (.A(G245P98gat), .Y(GB13gat) );
INVXL U_gB14 (.A(G552P152gat), .Y(GB14gat) );
INVXL U_gB15 (.A(G562P155gat), .Y(GB15gat) );
INVXL U_gB16 (.A(G559P154gat), .Y(GB16gat) );
INVXL U_gB17 (.A(G633P365gat), .Y(GB17gat) );
INVXL U_g3173P164_b (.A(G3173P164gat), .Y(G3173P164_bgat) );
AND2XL U_gB18 (.A(G136P62gat), .B(G3173P164_bgat), .Y(GB18gat) );
INVXL U_gB19 (.A(G844P657gat), .Y(GB19gat) );
INVXL U_gB20 (.A(G846P254gat), .Y(GB20gat) );
INVXL U_gB26 (.A(G549P151gat), .Y(GB26gat) );
INVXL U_g140P64_b (.A(G140P64gat), .Y(G140P64_bgat) );
INVXL U_g2822P361_b (.A(G2822P361gat), .Y(G2822P361_bgat) );
OR2XL U_gB27 (.A(G140P64_bgat), .B(G2822P361_bgat), .Y(GB27gat) );
INVXL U_gB28 (.A(G2822P361gat), .Y(GB28gat) );
INVXL U_gB34 (.A(G299P113gat), .Y(GB34gat) );
INVXL U_gB35 (.A(G635P1114gat), .Y(GB35gat) );
INVXL U_gB36 (.A(G703P1115gat), .Y(GB36gat) );
INVXL U_gB37 (.A(G716P1116gat), .Y(GB37gat) );
INVXL U_gB38 (.A(G819P1117gat), .Y(GB38gat) );
AND2XL U_gB39 (.A(G141P65gat), .B(G637P965gat), .Y(GB39gat) );
AND2XL U_gB40 (.A(G141P65gat), .B(G671P966gat), .Y(GB40gat) );
AND2XL U_gB41 (.A(G141P65gat), .B(G705P964gat), .Y(GB41gat) );
AND2XL U_gB42 (.A(G141P65gat), .B(G713P967gat), .Y(GB42gat) );
AND3XL U_gB43 (.A(G595P1463gat), .B(G596P1412gat), .C(G3328P916gat), .Y(GB43gat) );
INVXL U_g3350P1331_b (.A(G3350P1331gat), .Y(G3350P1331_bgat) );
AND3XL U_gB44 (.A(G607P1425gat), .B(G608P1440gat), .C(G3350P1331_bgat), .Y(GB44gat) );
AND2XL U_gB45 (.A(G1437P1530gat), .B(G1451P1551gat), .Y(GB45gat) );
AND2XL U_gB46 (.A(G1843P1630gat), .B(G1857P1608gat), .Y(GB46gat) );
AND2XL U_gB47 (.A(G2113P1632gat), .B(G2128P1619gat), .Y(GB47gat) );
AND2XL U_gB48 (.A(G1166P1522gat), .B(G1179P1552gat), .Y(GB48gat) );
INVXL U_g3532P1627_b (.A(G3532P1627gat), .Y(G3532P1627_bgat) );
INVXL U_g3531P1757_b (.A(G3531P1757gat), .Y(G3531P1757_bgat) );
OR2XL U_gB49 (.A(G3532P1627_bgat), .B(G3531P1757_bgat), .Y(GB49gat) );
INVXL U_g3967P1769_b (.A(G3967P1769gat), .Y(G3967P1769_bgat) );
INVXL U_g3966P1862_b (.A(G3966P1862gat), .Y(G3966P1862_bgat) );
OR2XL U_gB50 (.A(G3967P1769_bgat), .B(G3966P1862_bgat), .Y(GB50gat) );
OR2XL U_gB51 (.A(G589P1711gat), .B(G590P1806gat), .Y(GB51gat) );
OR2XL U_gB52 (.A(G616P1763gat), .B(G617P1849gat), .Y(GB52gat) );
OR2XL U_gB53 (.A(G619P1710gat), .B(G620P1800gat), .Y(GB53gat) );
OR2XL U_gB54 (.A(G627P1764gat), .B(G628P1853gat), .Y(GB54gat) );
INVXL U_gB55 (.A(G3848P1864gat), .Y(GB55gat) );
INVXL U_gB56 (.A(G3849P2024gat), .Y(GB56gat) );
INVXL U_gB57 (.A(G3790P2025gat), .Y(GB57gat) );
INVXL U_gB58 (.A(G1936P2105gat), .Y(GB58gat) );
OR4XL U_gB59 (.A(G718P1867gat), .B(G719P2030gat), .C(G720P848gat), .D(G721P646gat), .Y(GB59gat) );
INVXL U_gB60 (.A(G4082P2071gat), .Y(GB60gat) );
INVXL U_gB61 (.A(G3851P2063gat), .Y(GB61gat) );
INVXL U_gB62 (.A(G3850P2069gat), .Y(GB62gat) );
OR4XL U_gB63 (.A(G855P1866gat), .B(G856P2029gat), .C(G857P849gat), .D(G858P647gat), .Y(GB63gat) );
INVXL U_gB64 (.A(G4024P2068gat), .Y(GB64gat) );
INVXL U_gB65 (.A(G3793P2065gat), .Y(GB65gat) );
INVXL U_gB66 (.A(G3792P2066gat), .Y(GB66gat) );
INVXL U_gB67 (.A(G3791P2067gat), .Y(GB67gat) );
INVXL U_g3537P2019_b (.A(G3537P2019gat), .Y(G3537P2019_bgat) );
INVXL U_g3536P2059_b (.A(G3536P2059gat), .Y(G3536P2059_bgat) );
OR2XL U_gB68 (.A(G3537P2019_bgat), .B(G3536P2059_bgat), .Y(GB68gat) );
INVXL U_g3542P2023_b (.A(G3542P2023gat), .Y(G3542P2023_bgat) );
INVXL U_g3541P2062_b (.A(G3541P2062gat), .Y(G3541P2062_bgat) );
OR2XL U_gB69 (.A(G3542P2023_bgat), .B(G3541P2062_bgat), .Y(GB69gat) );
INVXL U_g1200P1934_b (.A(G1200P1934gat), .Y(G1200P1934_bgat) );
INVXL U_g1238P1953_b (.A(G1238P1953gat), .Y(G1238P1953_bgat) );
INVXL U_g1248P1959_b (.A(G1248P1959gat), .Y(G1248P1959_bgat) );
INVXL U_g1253P1960_b (.A(G1253P1960gat), .Y(G1253P1960_bgat) );
INVXL U_g1243P1961_b (.A(G1243P1961gat), .Y(G1243P1961_bgat) );
INVXL U_g1273P2005_b (.A(G1273P2005gat), .Y(G1273P2005_bgat) );
INVXL U_g1268P2050_b (.A(G1268P2050gat), .Y(G1268P2050_bgat) );
INVXL U_g1263P2111_b (.A(G1263P2111gat), .Y(G1263P2111_bgat) );
INVXL U_g1258P2112_b (.A(G1258P2112gat), .Y(G1258P2112_bgat) );
AND9XL U_gB70 (.A(G1200P1934_bgat), .B(G1238P1953_bgat), .C(G1248P1959_bgat), .D(G1253P1960_bgat), .E(G1243P1961_bgat), .F(G1273P2005_bgat), .G(G1268P2050_bgat), .H(G1263P2111_bgat), .I(G1258P2112_bgat), .Y(GB70gat) );
INVXL U_g1936P2105_b (.A(G1936P2105gat), .Y(G1936P2105_bgat) );
INVXL U_g1878P1647_b (.A(G1878P1647gat), .Y(G1878P1647_bgat) );
INVXL U_g1931P1914_b (.A(G1931P1914gat), .Y(G1931P1914_bgat) );
INVXL U_g1926P1937_b (.A(G1926P1937gat), .Y(G1926P1937_bgat) );
INVXL U_g1921P1939_b (.A(G1921P1939gat), .Y(G1921P1939_bgat) );
INVXL U_g1916P1940_b (.A(G1916P1940gat), .Y(G1916P1940_bgat) );
INVXL U_g1954P1997_b (.A(G1954P1997gat), .Y(G1954P1997_bgat) );
INVXL U_g1949P2040_b (.A(G1949P2040gat), .Y(G1949P2040_bgat) );
INVXL U_g1944P2104_b (.A(G1944P2104gat), .Y(G1944P2104_bgat) );
AND9XL U_gB71 (.A(G1936P2105_bgat), .B(G1878P1647_bgat), .C(G1931P1914_bgat), .D(G1926P1937_bgat), .E(G1921P1939_bgat), .F(G1916P1940_bgat), .G(G1954P1997_bgat), .H(G1949P2040_bgat), .I(G1944P2104_bgat), .Y(GB71gat) );
AND2XL U_gB72 (.A(G137P63gat), .B(G659P2121gat), .Y(GB72gat) );
AND2XL U_gB73 (.A(G137P63gat), .B(G691P2122gat), .Y(GB73gat) );
OR4XL U_gB74 (.A(G743P2082gat), .B(G744P2081gat), .C(G745P841gat), .D(G746P654gat), .Y(GB74gat) );
OR4XL U_gB75 (.A(G748P2086gat), .B(G749P2083gat), .C(G750P831gat), .D(G751P659gat), .Y(GB75gat) );
OR4XL U_gB76 (.A(G753P2087gat), .B(G754P2084gat), .C(G755P832gat), .D(G756P660gat), .Y(GB76gat) );
OR4XL U_gB77 (.A(G758P2031gat), .B(G759P2085gat), .C(G760P835gat), .D(G761P643gat), .Y(GB77gat) );
OR4XL U_gB78 (.A(G783P2074gat), .B(G784P2077gat), .C(G785P840gat), .D(G786P653gat), .Y(GB78gat) );
OR4XL U_gB79 (.A(G788P2075gat), .B(G789P2078gat), .C(G790P830gat), .D(G791P658gat), .Y(GB79gat) );
OR4XL U_gB80 (.A(G793P2076gat), .B(G794P2079gat), .C(G795P833gat), .D(G796P661gat), .Y(GB80gat) );
OR4XL U_gB81 (.A(G798P2028gat), .B(G799P2080gat), .C(G800P834gat), .D(G801P642gat), .Y(GB81gat) );
AND2XL U_gB82 (.A(G137P63gat), .B(G640P2170gat), .Y(GB82gat) );
AND2XL U_gB83 (.A(G137P63gat), .B(G662P2173gat), .Y(GB83gat) );
AND2XL U_gB84 (.A(G137P63gat), .B(G665P2174gat), .Y(GB84gat) );
AND2XL U_gB85 (.A(G137P63gat), .B(G668P2177gat), .Y(GB85gat) );
AND2XL U_gB86 (.A(G137P63gat), .B(G674P2171gat), .Y(GB86gat) );
AND2XL U_gB87 (.A(G137P63gat), .B(G694P2172gat), .Y(GB87gat) );
AND2XL U_gB88 (.A(G137P63gat), .B(G697P2175gat), .Y(GB88gat) );
AND2XL U_gB89 (.A(G137P63gat), .B(G700P2176gat), .Y(GB89gat) );
INVXL U_g4114P359_b (.A(G4114P359gat), .Y(G4114P359_bgat) );
AND2XL U_gB90 (.A(G817P2230gat), .B(G4114P359_bgat), .Y(GB90gat) );
OR2XL U_gB91 (.A(G811P2219gat), .B(G812P2205gat), .Y(GB91gat) );
INVXL U_gB92 (.A(G4086P2231gat), .Y(GB92gat) );
INVXL U_gB93 (.A(G4085P2232gat), .Y(GB93gat) );
INVXL U_gB94 (.A(G4084P2180gat), .Y(GB94gat) );
INVXL U_gB95 (.A(G4083P2130gat), .Y(GB95gat) );
AND3XL U_gB96 (.A(G245P98gat), .B(G852P255gat), .C(G853P2202gat), .Y(GB96gat) );
INVXL U_gB97 (.A(G4028P2234gat), .Y(GB97gat) );
INVXL U_gB98 (.A(G4027P2235gat), .Y(GB98gat) );
INVXL U_gB99 (.A(G4026P2185gat), .Y(GB99gat) );
INVXL U_gB100 (.A(G4025P2129gat), .Y(GB100gat) );
OR4XL U_gB101 (.A(G708P2243gat), .B(G709P2245gat), .C(G710P822gat), .D(G711P630gat), .Y(GB101gat) );
OR4XL U_gB102 (.A(G723P2249gat), .B(G724P2247gat), .C(G725P823gat), .D(G726P631gat), .Y(GB102gat) );
OR4XL U_gB103 (.A(G728P2250gat), .B(G729P2248gat), .C(G730P839gat), .D(G731P650gat), .Y(GB103gat) );
OR4XL U_gB104 (.A(G733P2197gat), .B(G734P2196gat), .C(G735P825gat), .D(G736P633gat), .Y(GB104gat) );
OR4XL U_gB105 (.A(G738P2141gat), .B(G739P2140gat), .C(G740P827gat), .D(G741P651gat), .Y(GB105gat) );
OR4XL U_gB106 (.A(G768P2244gat), .B(G769P2246gat), .C(G770P838gat), .D(G771P649gat), .Y(GB106gat) );
OR4XL U_gB107 (.A(G773P2194gat), .B(G774P2195gat), .C(G775P824gat), .D(G776P632gat), .Y(GB107gat) );
OR4XL U_gB108 (.A(G778P2138gat), .B(G779P2139gat), .C(G780P826gat), .D(G781P652gat), .Y(GB108gat) );
AND2XL U_gB109 (.A(G137P63gat), .B(G643P2221gat), .Y(GB109gat) );
AND2XL U_gB110 (.A(G137P63gat), .B(G646P2269gat), .Y(GB110gat) );
AND2XL U_gB111 (.A(G137P63gat), .B(G649P2292gat), .Y(GB111gat) );
AND2XL U_gB112 (.A(G137P63gat), .B(G652P2293gat), .Y(GB112gat) );
AND2XL U_gB113 (.A(G137P63gat), .B(G677P2220gat), .Y(GB113gat) );
AND2XL U_gB114 (.A(G137P63gat), .B(G680P2270gat), .Y(GB114gat) );
AND2XL U_gB115 (.A(G137P63gat), .B(G683P2291gat), .Y(GB115gat) );
AND2XL U_gB116 (.A(G137P63gat), .B(G686P2294gat), .Y(GB116gat) );
OR4XL U_gB117 (.A(G839P2241gat), .B(G840P2451gat), .C(G841P813gat), .D(G842P368gat), .Y(GB117gat) );
OR4XL U_gB118 (.A(G878P2242gat), .B(G879P2452gat), .C(G880P815gat), .D(G881P370gat), .Y(GB118gat) );
OR4XL U_gB119 (.A(G763P2472gat), .B(G764P2471gat), .C(G765P847gat), .D(G766P644gat), .Y(GB119gat) );
OR4XL U_gB120 (.A(G803P2469gat), .B(G804P2470gat), .C(G805P846gat), .D(G806P645gat), .Y(GB120gat) );
INVXL U_gB121 (.A(G657P2481gat), .Y(GB121gat) );
INVXL U_gB122 (.A(G689P2482gat), .Y(GB122gat) );
INVXL U_g1P0_b (.A(G1P0gat), .Y(G1P0_bgat) );
INVXL U_g373P133_b (.A(G373P133gat), .Y(G373P133_bgat) );
OR2XL U_g633P365 (.A(G1P0_bgat), .B(G373P133_bgat), .Y(G633P365gat) );
INVXL U_g2824P163_b (.A(G2824P163gat), .Y(G2824P163_bgat) );
AND2XL U_g844P657 (.A(G27P10gat), .B(G2824P163_bgat), .Y(G844P657gat) );
AND2XL U_g846P254 (.A(G386P135gat), .B(G556P153gat), .Y(G846P254gat) );
AND2XL U_g2822P361 (.A(G27P10gat), .B(G31P11gat), .Y(G2822P361gat) );
AND2XL U_g635P1114 (.A(G3176P362gat), .B(G3197P953gat), .Y(G635P1114gat) );
AND2XL U_g703P1115 (.A(G3176P362gat), .B(G3200P952gat), .Y(G703P1115gat) );
AND2XL U_g716P1116 (.A(G3176P362gat), .B(G3203P951gat), .Y(G716P1116gat) );
AND2XL U_g819P1117 (.A(G3176P362gat), .B(G3194P954gat), .Y(G819P1117gat) );
OR4XL U_g637P965 (.A(G2881P678gat), .B(G2880P684gat), .C(G2879P960gat), .D(G2878P961gat), .Y(G637P965gat) );
OR4XL U_g671P966 (.A(G2877P679gat), .B(G2876P683gat), .C(G2875P956gat), .D(G2874P959gat), .Y(G671P966gat) );
OR4XL U_g705P964 (.A(G2869P677gat), .B(G2868P681gat), .C(G2866P958gat), .D(G2867P962gat), .Y(G705P964gat) );
OR4XL U_g713P967 (.A(G2873P680gat), .B(G2872P682gat), .C(G2870P955gat), .D(G2871P957gat), .Y(G713P967gat) );
INVXL U_g2933P933_b (.A(G2933P933gat), .Y(G2933P933_bgat) );
INVXL U_g2942P1137_b (.A(G2942P1137gat), .Y(G2942P1137_bgat) );
INVXL U_g2939P1144_b (.A(G2939P1144gat), .Y(G2939P1144_bgat) );
AND4XL U_g595P1463 (.A(G2908P930gat), .B(G2933P933_bgat), .C(G2942P1137_bgat), .D(G2939P1144_bgat), .Y(G595P1463gat) );
INVXL U_g3015P863_b (.A(G3015P863gat), .Y(G3015P863_bgat) );
INVXL U_g3021P1123_b (.A(G3021P1123gat), .Y(G3021P1123_bgat) );
INVXL U_g3018P1126_b (.A(G3018P1126gat), .Y(G3018P1126_bgat) );
INVXL U_g3012P1132_b (.A(G3012P1132gat), .Y(G3012P1132_bgat) );
AND4XL U_g596P1412 (.A(G3015P863_bgat), .B(G3021P1123_bgat), .C(G3018P1126_bgat), .D(G3012P1132_bgat), .Y(G596P1412gat) );
INVXL U_g2615P1155_b (.A(G2615P1155gat), .Y(G2615P1155_bgat) );
INVXL U_g2611P1159_b (.A(G2611P1159gat), .Y(G2611P1159_bgat) );
INVXL U_g2623P1167_b (.A(G2623P1167gat), .Y(G2623P1167_bgat) );
INVXL U_g2619P1171_b (.A(G2619P1171gat), .Y(G2619P1171_bgat) );
AND4XL U_g607P1425 (.A(G2615P1155_bgat), .B(G2611P1159_bgat), .C(G2623P1167_bgat), .D(G2619P1171_bgat), .Y(G607P1425gat) );
INVXL U_g2713P1178_b (.A(G2713P1178gat), .Y(G2713P1178_bgat) );
INVXL U_g2709P1183_b (.A(G2709P1183gat), .Y(G2709P1183_bgat) );
INVXL U_g2705P1186_b (.A(G2705P1186gat), .Y(G2705P1186_bgat) );
INVXL U_g2717P1191_b (.A(G2717P1191gat), .Y(G2717P1191_bgat) );
AND4XL U_g608P1440 (.A(G2713P1178_bgat), .B(G2709P1183_bgat), .C(G2705P1186_bgat), .D(G2717P1191_bgat), .Y(G608P1440gat) );
AND4XL U_g1437P1530 (.A(G1307P1427gat), .B(G1289P1428gat), .C(G1278P1433gat), .D(G1422P1439gat), .Y(G1437P1530gat) );
AND5XL U_g1451P1551 (.A(G1332P1435gat), .B(G1390P1443gat), .C(G1365P1445gat), .D(G1344P1449gat), .E(G1430P1451gat), .Y(G1451P1551gat) );
INVXL U_g3165P927_b (.A(G3165P927gat), .Y(G3165P927_bgat) );
INVXL U_g3167P931_b (.A(G3167P931gat), .Y(G3167P931_bgat) );
AND4XL U_g1843P1630 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G1758P1420gat), .D(G1730P1422gat), .Y(G1843P1630gat) );
INVXL U_g3137P914_b (.A(G3137P914gat), .Y(G3137P914_bgat) );
AND5XL U_g1857P1608 (.A(G3137P914_bgat), .B(G1778P1307gat), .C(G1812P1404gat), .D(G1794P1406gat), .E(G1767P1417gat), .Y(G1857P1608gat) );
AND4XL U_g2113P1632 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G2099P1419gat), .D(G1984P1423gat), .Y(G2113P1632gat) );
AND5XL U_g2128P1619 (.A(G3137P914_bgat), .B(G2021P1306gat), .C(G2067P1403gat), .D(G2042P1408gat), .E(G2009P1416gat), .Y(G2128P1619gat) );
AND4XL U_g1166P1522 (.A(G1052P1426gat), .B(G1034P1429gat), .C(G1023P1432gat), .D(G1080P1438gat), .Y(G1166P1522gat) );
AND5XL U_g1179P1552 (.A(G1089P1436gat), .B(G1134P1442gat), .C(G1116P1446gat), .D(G1100P1448gat), .E(G1152P1452gat), .Y(G1179P1552gat) );
OR4XL U_g589P1711 (.A(G1286P1007gat), .B(G1440P1534gat), .C(G1439P1539gat), .D(G1441P1563gat), .Y(G589P1711gat) );
AND2XL U_g590P1806 (.A(G1437P1530gat), .B(G1458P1719gat), .Y(G590P1806gat) );
OR4XL U_g616P1763 (.A(G3167P931gat), .B(G1846P1147gat), .C(G1845P1226gat), .D(G1847P1509gat), .Y(G616P1763gat) );
AND2XL U_g617P1849 (.A(G1843P1630gat), .B(G1863P1675gat), .Y(G617P1849gat) );
OR4XL U_g619P1710 (.A(G1031P1006gat), .B(G1169P1525gat), .C(G1168P1542gat), .D(G1170P1555gat), .Y(G619P1710gat) );
AND2XL U_g620P1800 (.A(G1166P1522gat), .B(G1185P1721gat), .Y(G620P1800gat) );
OR4XL U_g627P1764 (.A(G3167P931gat), .B(G2116P1152gat), .C(G2115P1229gat), .D(G2117P1504gat), .Y(G627P1764gat) );
AND2XL U_g628P1853 (.A(G2113P1632gat), .B(G2135P1673gat), .Y(G628P1853gat) );
OR3XL U_g3848P1864 (.A(G3838P804gat), .B(G3836P1120gat), .C(G3837P1653gat), .Y(G3848P1864gat) );
OR3XL U_g3849P2024 (.A(G3841P806gat), .B(G3839P1291gat), .C(G3840P1935gat), .Y(G3849P2024gat) );
OR3XL U_g3790P2025 (.A(G3780P816gat), .B(G3778P1293gat), .C(G3779P1936gat), .Y(G3790P2025gat) );
OR2XL U_g1936P2105 (.A(G1935P1994gat), .B(G1934P2039gat), .Y(G1936P2105gat) );
INVXL U_g4087P171_b (.A(G4087P171gat), .Y(G4087P171_bgat) );
INVXL U_g4088P172_b (.A(G4088P172gat), .Y(G4088P172_bgat) );
AND3XL U_g718P1867 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G3848P1864gat), .Y(G718P1867gat) );
AND3XL U_g719P2030 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G3790P2025gat), .Y(G719P2030gat) );
AND3XL U_g720P848 (.A(G11P2gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G720P848gat) );
AND3XL U_g721P646 (.A(G61P21gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G721P646gat) );
OR3XL U_g4082P2071 (.A(G4069P837gat), .B(G4067P1284gat), .C(G4068P1980gat), .Y(G4082P2071gat) );
OR3XL U_g3851P2063 (.A(G3847P805gat), .B(G3845P963gat), .C(G3846P1982gat), .Y(G3851P2063gat) );
OR3XL U_g3850P2069 (.A(G3844P814gat), .B(G3842P1292gat), .C(G3843P1983gat), .Y(G3850P2069gat) );
INVXL U_g4089P173_b (.A(G4089P173gat), .Y(G4089P173_bgat) );
INVXL U_g4090P174_b (.A(G4090P174gat), .Y(G4090P174_bgat) );
AND3XL U_g855P1866 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G3848P1864gat), .Y(G855P1866gat) );
AND3XL U_g856P2029 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G3790P2025gat), .Y(G856P2029gat) );
AND3XL U_g857P849 (.A(G11P2gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G857P849gat) );
AND3XL U_g858P647 (.A(G61P21gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G858P647gat) );
OR3XL U_g4024P2068 (.A(G4011P811gat), .B(G4009P1287gat), .C(G4010P1981gat), .Y(G4024P2068gat) );
OR3XL U_g3793P2065 (.A(G3789P807gat), .B(G3787P1296gat), .C(G3788P1984gat), .Y(G3793P2065gat) );
OR3XL U_g3792P2066 (.A(G3786P808gat), .B(G3784P1295gat), .C(G3785P1985gat), .Y(G3792P2066gat) );
OR3XL U_g3791P2067 (.A(G3783P809gat), .B(G3781P1294gat), .C(G3782P1986gat), .Y(G3791P2067gat) );
OR4XL U_g659P2121 (.A(G1668P599gat), .B(G1667P797gat), .C(G1664P1870gat), .D(G1666P2035gat), .Y(G659P2121gat) );
OR4XL U_g691P2122 (.A(G2339P600gat), .B(G2338P796gat), .C(G2335P1869gat), .D(G2337P2033gat), .Y(G691P2122gat) );
AND3XL U_g743P2082 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G4082P2071gat), .Y(G743P2082gat) );
AND3XL U_g744P2081 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G4024P2068gat), .Y(G744P2081gat) );
AND3XL U_g745P841 (.A(G43P15gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G745P841gat) );
AND3XL U_g746P654 (.A(G37P13gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G746P654gat) );
AND3XL U_g748P2086 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G3851P2063gat), .Y(G748P2086gat) );
AND3XL U_g749P2083 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G3793P2065gat), .Y(G749P2083gat) );
AND3XL U_g750P831 (.A(G76P26gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G750P831gat) );
AND3XL U_g751P659 (.A(G20P5gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G751P659gat) );
AND3XL U_g753P2087 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G3850P2069gat), .Y(G753P2087gat) );
AND3XL U_g754P2084 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G3792P2066gat), .Y(G754P2084gat) );
AND3XL U_g755P832 (.A(G73P25gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G755P832gat) );
AND3XL U_g756P660 (.A(G17P4gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G756P660gat) );
AND3XL U_g758P2031 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G3849P2024gat), .Y(G758P2031gat) );
AND3XL U_g759P2085 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G3791P2067gat), .Y(G759P2085gat) );
AND3XL U_g760P835 (.A(G67P23gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G760P835gat) );
AND3XL U_g761P643 (.A(G70P24gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G761P643gat) );
AND3XL U_g783P2074 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G4082P2071gat), .Y(G783P2074gat) );
AND3XL U_g784P2077 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G4024P2068gat), .Y(G784P2077gat) );
AND3XL U_g785P840 (.A(G43P15gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G785P840gat) );
AND3XL U_g786P653 (.A(G37P13gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G786P653gat) );
AND3XL U_g788P2075 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G3851P2063gat), .Y(G788P2075gat) );
AND3XL U_g789P2078 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G3793P2065gat), .Y(G789P2078gat) );
AND3XL U_g790P830 (.A(G76P26gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G790P830gat) );
AND3XL U_g791P658 (.A(G20P5gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G791P658gat) );
AND3XL U_g793P2076 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G3850P2069gat), .Y(G793P2076gat) );
AND3XL U_g794P2079 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G3792P2066gat), .Y(G794P2079gat) );
AND3XL U_g795P833 (.A(G73P25gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G795P833gat) );
AND3XL U_g796P661 (.A(G17P4gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G796P661gat) );
AND3XL U_g798P2028 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G3849P2024gat), .Y(G798P2028gat) );
AND3XL U_g799P2080 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G3791P2067gat), .Y(G799P2080gat) );
AND3XL U_g800P834 (.A(G67P23gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G800P834gat) );
AND3XL U_g801P642 (.A(G70P24gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G801P642gat) );
OR4XL U_g640P2170 (.A(G1580P605gat), .B(G1579P787gat), .C(G1576P2097gat), .D(G1578P2101gat), .Y(G640P2170gat) );
OR4XL U_g662P2173 (.A(G1674P614gat), .B(G1673P794gat), .C(G1670P2034gat), .D(G1672P2100gat), .Y(G662P2173gat) );
OR4XL U_g665P2174 (.A(G1680P615gat), .B(G1679P801gat), .C(G1676P2095gat), .D(G1678P2099gat), .Y(G665P2174gat) );
OR4XL U_g668P2177 (.A(G1686P618gat), .B(G1685P802gat), .C(G1682P2096gat), .D(G1684P2098gat), .Y(G668P2177gat) );
OR4XL U_g674P2171 (.A(G2254P606gat), .B(G2253P786gat), .C(G2250P2090gat), .D(G2252P2094gat), .Y(G674P2171gat) );
OR4XL U_g694P2172 (.A(G2345P613gat), .B(G2344P795gat), .C(G2341P2032gat), .D(G2343P2093gat), .Y(G694P2172gat) );
OR4XL U_g697P2175 (.A(G2351P616gat), .B(G2350P800gat), .C(G2347P2088gat), .D(G2349P2092gat), .Y(G697P2175gat) );
OR4XL U_g700P2176 (.A(G2357P617gat), .B(G2356P803gat), .C(G2353P2089gat), .D(G2355P2091gat), .Y(G700P2176gat) );
OR4XL U_g817P2230 (.A(G3734P629gat), .B(G3731P1121gat), .C(G3733P1868gat), .D(G3735P2142gat), .Y(G817P2230gat) );
AND2XL U_g811P2219 (.A(G4113P1859gat), .B(G4096P2167gat), .Y(G811P2219gat) );
AND2XL U_g812P2205 (.A(G1936P2105gat), .B(G4096P2167gat), .Y(G812P2205gat) );
OR3XL U_g4086P2231 (.A(G4081P810gat), .B(G4079P1119gat), .C(G4080P2134gat), .Y(G4086P2231gat) );
OR3XL U_g4085P2232 (.A(G4078P812gat), .B(G4076P1118gat), .C(G4077P2135gat), .Y(G4085P2232gat) );
OR3XL U_g4084P2180 (.A(G4075P817gat), .B(G4073P1286gat), .C(G4074P2072gat), .Y(G4084P2180gat) );
OR3XL U_g4083P2130 (.A(G4072P821gat), .B(G4070P1285gat), .C(G4071P2026gat), .Y(G4083P2130gat) );
AND4XL U_g852P255 (.A(G386P135gat), .B(G552P152gat), .C(G556P153gat), .D(G559P154gat), .Y(G852P255gat) );
INVXL U_gB49_b (.A(GB49gat), .Y(GB49_bgat) );
INVXL U_gB50_b (.A(GB50gat), .Y(GB50_bgat) );
INVXL U_gB68_b (.A(GB68gat), .Y(GB68_bgat) );
INVXL U_gB69_b (.A(GB69gat), .Y(GB69_bgat) );
AND5XL U_g853P2202 (.A(G562P155gat), .B(GB49_bgat), .C(GB50_bgat), .D(GB68_bgat), .E(GB69_bgat), .Y(G853P2202gat) );
OR3XL U_g4028P2234 (.A(G4023P818gat), .B(G4021P1401gat), .C(G4022P2136gat), .Y(G4028P2234gat) );
OR3XL U_g4027P2235 (.A(G4020P819gat), .B(G4018P1290gat), .C(G4019P2137gat), .Y(G4027P2235gat) );
OR3XL U_g4026P2185 (.A(G4017P836gat), .B(G4015P1289gat), .C(G4016P2073gat), .Y(G4026P2185gat) );
OR3XL U_g4025P2129 (.A(G4014P820gat), .B(G4012P1288gat), .C(G4013P2027gat), .Y(G4025P2129gat) );
AND3XL U_g708P2243 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G4086P2231gat), .Y(G708P2243gat) );
AND3XL U_g709P2245 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G4028P2234gat), .Y(G709P2245gat) );
AND3XL U_g710P822 (.A(G109P41gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G710P822gat) );
AND3XL U_g711P630 (.A(G106P40gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G711P630gat) );
AND3XL U_g723P2249 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G4086P2231gat), .Y(G723P2249gat) );
AND3XL U_g724P2247 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G4028P2234gat), .Y(G724P2247gat) );
AND3XL U_g725P823 (.A(G109P41gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G725P823gat) );
AND3XL U_g726P631 (.A(G106P40gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G726P631gat) );
AND3XL U_g728P2250 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G4085P2232gat), .Y(G728P2250gat) );
AND3XL U_g729P2248 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G4027P2235gat), .Y(G729P2248gat) );
AND3XL U_g730P839 (.A(G46P16gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G730P839gat) );
AND3XL U_g731P650 (.A(G49P17gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G731P650gat) );
AND3XL U_g733P2197 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G4084P2180gat), .Y(G733P2197gat) );
AND3XL U_g734P2196 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G4026P2185gat), .Y(G734P2196gat) );
AND3XL U_g735P825 (.A(G100P38gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G735P825gat) );
AND3XL U_g736P633 (.A(G103P39gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G736P633gat) );
AND3XL U_g738P2141 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G4083P2130gat), .Y(G738P2141gat) );
AND3XL U_g739P2140 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G4025P2129gat), .Y(G739P2140gat) );
AND3XL U_g740P827 (.A(G91P35gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G740P827gat) );
AND3XL U_g741P651 (.A(G40P14gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G741P651gat) );
AND3XL U_g768P2244 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G4085P2232gat), .Y(G768P2244gat) );
AND3XL U_g769P2246 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G4027P2235gat), .Y(G769P2246gat) );
AND3XL U_g770P838 (.A(G46P16gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G770P838gat) );
AND3XL U_g771P649 (.A(G49P17gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G771P649gat) );
AND3XL U_g773P2194 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G4084P2180gat), .Y(G773P2194gat) );
AND3XL U_g774P2195 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G4026P2185gat), .Y(G774P2195gat) );
AND3XL U_g775P824 (.A(G100P38gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G775P824gat) );
AND3XL U_g776P632 (.A(G103P39gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G776P632gat) );
AND3XL U_g778P2138 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G4083P2130gat), .Y(G778P2138gat) );
AND3XL U_g779P2139 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G4025P2129gat), .Y(G779P2139gat) );
AND3XL U_g780P826 (.A(G91P35gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G780P826gat) );
AND3XL U_g781P652 (.A(G40P14gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G781P652gat) );
OR4XL U_g643P2221 (.A(G1586P604gat), .B(G1585P785gat), .C(G1582P2145gat), .D(G1584P2146gat), .Y(G643P2221gat) );
OR4XL U_g646P2269 (.A(G1592P607gat), .B(G1591P789gat), .C(G1588P2200gat), .D(G1590P2201gat), .Y(G646P2269gat) );
OR4XL U_g649P2292 (.A(G1598P610gat), .B(G1597P791gat), .C(G1594P2255gat), .D(G1596P2258gat), .Y(G649P2292gat) );
OR4XL U_g652P2293 (.A(G1604P611gat), .B(G1603P793gat), .C(G1600P2256gat), .D(G1602P2257gat), .Y(G652P2293gat) );
OR4XL U_g677P2220 (.A(G2260P603gat), .B(G2259P784gat), .C(G2256P2143gat), .D(G2258P2144gat), .Y(G677P2220gat) );
OR4XL U_g680P2270 (.A(G2266P608gat), .B(G2265P788gat), .C(G2262P2198gat), .D(G2264P2199gat), .Y(G680P2270gat) );
OR4XL U_g683P2291 (.A(G2272P609gat), .B(G2271P790gat), .C(G2268P2251gat), .D(G2270P2254gat), .Y(G683P2291gat) );
OR4XL U_g686P2294 (.A(G2278P612gat), .B(G2277P792gat), .C(G2274P2252gat), .D(G2276P2253gat), .Y(G686P2294gat) );
INVXL U_g4091P175_b (.A(G4091P175gat), .Y(G4091P175_bgat) );
INVXL U_g4092P176_b (.A(G4092P176gat), .Y(G4092P176_bgat) );
INVXL U_g3965P2153_b (.A(G3965P2153gat), .Y(G3965P2153_bgat) );
AND3XL U_g839P2241 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3965P2153_bgat), .Y(G839P2241gat) );
AND3XL U_g840P2451 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G2198P2449gat), .Y(G840P2451gat) );
AND3XL U_g841P813 (.A(G120P50gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G841P813gat) );
AND2XL U_g842P368 (.A(G4091P175gat), .B(G4092P176gat), .Y(G842P368gat) );
INVXL U_g3962P2154_b (.A(G3962P2154gat), .Y(G3962P2154_bgat) );
AND3XL U_g878P2242 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3962P2154_bgat), .Y(G878P2242gat) );
AND3XL U_g879P2452 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1521P2450gat), .Y(G879P2452gat) );
AND3XL U_g880P815 (.A(G118P48gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G880P815gat) );
AND2XL U_g881P370 (.A(G4091P175gat), .B(G4092P176gat), .Y(G881P370gat) );
AND3XL U_g763P2472 (.A(G4087P171_bgat), .B(G4088P172_bgat), .C(G3656P2467gat), .Y(G763P2472gat) );
AND3XL U_g764P2471 (.A(G4087P171_bgat), .B(G4088P172gat), .C(G3655P2465gat), .Y(G764P2471gat) );
AND3XL U_g765P847 (.A(G14P3gat), .B(G4087P171gat), .C(G4088P172_bgat), .Y(G765P847gat) );
AND3XL U_g766P644 (.A(G64P22gat), .B(G4087P171gat), .C(G4088P172gat), .Y(G766P644gat) );
AND3XL U_g803P2469 (.A(G4089P173_bgat), .B(G4090P174_bgat), .C(G3656P2467gat), .Y(G803P2469gat) );
AND3XL U_g804P2470 (.A(G4089P173gat), .B(G4090P174_bgat), .C(G3655P2465gat), .Y(G804P2470gat) );
AND3XL U_g805P846 (.A(G14P3gat), .B(G4089P173_bgat), .C(G4090P174gat), .Y(G805P846gat) );
AND3XL U_g806P645 (.A(G64P22gat), .B(G4089P173gat), .C(G4090P174gat), .Y(G806P645gat) );
AND2XL U_g657P2481 (.A(G137P63gat), .B(G1662P2477gat), .Y(G657P2481gat) );
AND2XL U_g689P2482 (.A(G137P63gat), .B(G2333P2478gat), .Y(G689P2482gat) );
AND2XL U_g4114P359 (.A(G135P61gat), .B(G4115P177gat), .Y(G4114P359gat) );
AND2XL U_g3176P362 (.A(G27P10gat), .B(G31P11gat), .Y(G3176P362gat) );
INVXL U_g3546P165_b (.A(G3546P165gat), .Y(G3546P165_bgat) );
AND2XL U_g2590P386 (.A(G210P89gat), .B(G3546P165_bgat), .Y(G2590P386gat) );
AND2XL U_g2595P387 (.A(G218P91gat), .B(G3546P165_bgat), .Y(G2595P387gat) );
AND2XL U_g2600P388 (.A(G226P93gat), .B(G3546P165_bgat), .Y(G2600P388gat) );
AND2XL U_g2605P389 (.A(G234P95gat), .B(G3546P165_bgat), .Y(G2605P389gat) );
AND2XL U_g2684P390 (.A(G257P102gat), .B(G3546P165_bgat), .Y(G2684P390gat) );
AND2XL U_g2689P391 (.A(G265P104gat), .B(G3546P165_bgat), .Y(G2689P391gat) );
AND2XL U_g2694P392 (.A(G273P106gat), .B(G3546P165_bgat), .Y(G2694P392gat) );
AND2XL U_g2699P393 (.A(G281P108gat), .B(G3546P165_bgat), .Y(G2699P393gat) );
AND2XL U_g2994P394 (.A(G324P120gat), .B(G3546P165_bgat), .Y(G2994P394gat) );
AND2XL U_g3001P395 (.A(G341P125gat), .B(G3546P165_bgat), .Y(G3001P395gat) );
AND2XL U_g3006P396 (.A(G351P127gat), .B(G3546P165_bgat), .Y(G3006P396gat) );
AND3XL U_g3238P409 (.A(G248P99gat), .B(G351P127gat), .C(G534P149gat), .Y(G3238P409gat) );
INVXL U_g3552P168_b (.A(G3552P168gat), .Y(G3552P168_bgat) );
AND3XL U_g2988P410 (.A(G351P127gat), .B(G534P149gat), .C(G3552P168_bgat), .Y(G2988P410gat) );
AND3XL U_g2982P413 (.A(G341P125gat), .B(G523P148gat), .C(G3552P168_bgat), .Y(G2982P413gat) );
AND3XL U_g3234P414 (.A(G248P99gat), .B(G341P125gat), .C(G523P148gat), .Y(G3234P414gat) );
OR2XL U_g3247P417 (.A(G242P97gat), .B(G514P147gat), .Y(G3247P417gat) );
AND2XL U_g3232P418 (.A(G248P99gat), .B(G514P147gat), .Y(G3232P418gat) );
OR2XL U_g2999P419 (.A(G514P147gat), .B(G3546P165_bgat), .Y(G2999P419gat) );
AND2XL U_g2979P420 (.A(G514P147gat), .B(G3552P168_bgat), .Y(G2979P420gat) );
AND3XL U_g2973P423 (.A(G324P120gat), .B(G503P146gat), .C(G3552P168_bgat), .Y(G2973P423gat) );
AND3XL U_g3228P424 (.A(G248P99gat), .B(G324P120gat), .C(G503P146gat), .Y(G3228P424gat) );
AND3XL U_g3287P427 (.A(G248P99gat), .B(G316P118gat), .C(G490P145gat), .Y(G3287P427gat) );
AND3XL U_g2913P428 (.A(G248P99gat), .B(G316P118gat), .C(G490P145gat), .Y(G2913P428gat) );
AND3XL U_g2909P431 (.A(G248P99gat), .B(G308P116gat), .C(G479P144gat), .Y(G2909P431gat) );
AND3XL U_g3283P432 (.A(G248P99gat), .B(G308P116gat), .C(G479P144gat), .Y(G3283P432gat) );
AND3XL U_g3390P435 (.A(G218P91gat), .B(G248P99gat), .C(G468P143gat), .Y(G3390P435gat) );
AND3XL U_g2572P436 (.A(G218P91gat), .B(G468P143gat), .C(G3552P168_bgat), .Y(G2572P436gat) );
AND3XL U_g3386P439 (.A(G210P89gat), .B(G248P99gat), .C(G457P142gat), .Y(G3386P439gat) );
AND3XL U_g2566P440 (.A(G210P89gat), .B(G457P142gat), .C(G3552P168_bgat), .Y(G2566P440gat) );
AND3XL U_g3398P445 (.A(G234P95gat), .B(G248P99gat), .C(G435P140gat), .Y(G3398P445gat) );
AND3XL U_g2584P446 (.A(G234P95gat), .B(G435P140gat), .C(G3552P168_bgat), .Y(G2584P446gat) );
AND3XL U_g3394P449 (.A(G226P93gat), .B(G248P99gat), .C(G422P139gat), .Y(G3394P449gat) );
AND3XL U_g2578P450 (.A(G226P93gat), .B(G422P139gat), .C(G3552P168_bgat), .Y(G2578P450gat) );
AND3XL U_g2672P453 (.A(G273P106gat), .B(G411P138gat), .C(G3552P168_bgat), .Y(G2672P453gat) );
AND3XL U_g3064P454 (.A(G248P99gat), .B(G273P106gat), .C(G411P138gat), .Y(G3064P454gat) );
AND3XL U_g3060P457 (.A(G248P99gat), .B(G265P104gat), .C(G400P137gat), .Y(G3060P457gat) );
AND3XL U_g2666P458 (.A(G265P104gat), .B(G400P137gat), .C(G3552P168_bgat), .Y(G2666P458gat) );
AND3XL U_g2660P461 (.A(G257P102gat), .B(G389P136gat), .C(G3552P168_bgat), .Y(G2660P461gat) );
AND3XL U_g3056P462 (.A(G248P99gat), .B(G257P102gat), .C(G389P136gat), .Y(G3056P462gat) );
AND3XL U_g3068P466 (.A(G248P99gat), .B(G281P108gat), .C(G374P134gat), .Y(G3068P466gat) );
AND3XL U_g2678P467 (.A(G281P108gat), .B(G374P134gat), .C(G3552P168_bgat), .Y(G2678P467gat) );
AND2XL U_g3119P470 (.A(G332P122gat), .B(G372P132gat), .Y(G3119P470gat) );
AND2XL U_g3121P472 (.A(G332P122gat), .B(G366P130gat), .Y(G3121P472gat) );
AND2XL U_g3333P473 (.A(G248P99gat), .B(G361P129gat), .Y(G3333P473gat) );
AND2XL U_g3326P475 (.A(G248P99gat), .B(G361P129gat), .Y(G3326P475gat) );
AND2XL U_g3123P478 (.A(G332P122gat), .B(G358P128gat), .Y(G3123P478gat) );
AND2XL U_g3253P480 (.A(G242P97gat), .B(G351P127gat), .Y(G3253P480gat) );
AND2XL U_g3125P485 (.A(G332P122gat), .B(G348P126gat), .Y(G3125P485gat) );
AND2XL U_g3249P486 (.A(G242P97gat), .B(G341P125gat), .Y(G3249P486gat) );
AND2XL U_g3126P492 (.A(G332P122gat), .B(G338P124gat), .Y(G3126P492gat) );
AND2XL U_g3128P497 (.A(G331P121gat), .B(G332P122gat), .Y(G3128P497gat) );
AND2XL U_g3243P498 (.A(G242P97gat), .B(G324P120gat), .Y(G3243P498gat) );
AND2XL U_g3130P505 (.A(G323P119gat), .B(G332P122gat), .Y(G3130P505gat) );
AND2XL U_g3299P507 (.A(G242P97gat), .B(G316P118gat), .Y(G3299P507gat) );
AND2XL U_g2927P510 (.A(G242P97gat), .B(G316P118gat), .Y(G2927P510gat) );
AND2XL U_g3132P513 (.A(G315P117gat), .B(G332P122gat), .Y(G3132P513gat) );
AND2XL U_g3295P515 (.A(G242P97gat), .B(G308P116gat), .Y(G3295P515gat) );
AND2XL U_g2922P518 (.A(G242P97gat), .B(G308P116gat), .Y(G2922P518gat) );
AND2XL U_g3134P521 (.A(G307P115gat), .B(G332P122gat), .Y(G3134P521gat) );
AND2XL U_g3280P522 (.A(G248P99gat), .B(G302P114gat), .Y(G3280P522gat) );
AND2XL U_g2906P525 (.A(G248P99gat), .B(G302P114gat), .Y(G2906P525gat) );
AND2XL U_g3136P529 (.A(G299P113gat), .B(G332P122gat), .Y(G3136P529gat) );
AND2XL U_g3292P531 (.A(G242P97gat), .B(G293P112gat), .Y(G3292P531gat) );
AND2XL U_g2918P533 (.A(G242P97gat), .B(G293P112gat), .Y(G2918P533gat) );
AND2XL U_g2748P535 (.A(G292P111gat), .B(G335P123gat), .Y(G2748P535gat) );
AND2XL U_g2750P537 (.A(G288P109gat), .B(G335P123gat), .Y(G2750P537gat) );
AND2XL U_g3088P539 (.A(G242P97gat), .B(G281P108gat), .Y(G3088P539gat) );
AND2XL U_g2752P544 (.A(G280P107gat), .B(G335P123gat), .Y(G2752P544gat) );
AND2XL U_g3083P545 (.A(G242P97gat), .B(G273P106gat), .Y(G3083P545gat) );
AND2XL U_g2754P551 (.A(G272P105gat), .B(G335P123gat), .Y(G2754P551gat) );
AND2XL U_g3078P553 (.A(G242P97gat), .B(G265P104gat), .Y(G3078P553gat) );
AND2XL U_g2756P558 (.A(G264P103gat), .B(G335P123gat), .Y(G2756P558gat) );
AND2XL U_g3073P560 (.A(G242P97gat), .B(G257P102gat), .Y(G3073P560gat) );
AND2XL U_g3403P565 (.A(G210P89gat), .B(G242P97gat), .Y(G3403P565gat) );
AND2XL U_g3408P566 (.A(G218P91gat), .B(G242P97gat), .Y(G3408P566gat) );
AND2XL U_g3413P567 (.A(G226P93gat), .B(G242P97gat), .Y(G3413P567gat) );
AND2XL U_g3418P568 (.A(G234P95gat), .B(G242P97gat), .Y(G3418P568gat) );
AND2XL U_g2758P569 (.A(G241P96gat), .B(G335P123gat), .Y(G2758P569gat) );
AND2XL U_g2760P575 (.A(G233P94gat), .B(G335P123gat), .Y(G2760P575gat) );
AND2XL U_g2762P581 (.A(G225P92gat), .B(G335P123gat), .Y(G2762P581gat) );
AND2XL U_g2764P587 (.A(G217P90gat), .B(G335P123gat), .Y(G2764P587gat) );
AND2XL U_g2766P593 (.A(G209P88gat), .B(G335P123gat), .Y(G2766P593gat) );
AND3XL U_g1668P599 (.A(G185P80gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1668P599gat) );
AND3XL U_g2339P600 (.A(G185P80gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2339P600gat) );
AND3XL U_g1661P601 (.A(G179P78gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1661P601gat) );
AND3XL U_g2332P602 (.A(G179P78gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2332P602gat) );
AND3XL U_g2260P603 (.A(G173P76gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2260P603gat) );
AND3XL U_g1586P604 (.A(G173P76gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1586P604gat) );
AND3XL U_g1580P605 (.A(G170P75gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1580P605gat) );
AND3XL U_g2254P606 (.A(G170P75gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2254P606gat) );
AND3XL U_g1592P607 (.A(G167P74gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1592P607gat) );
AND3XL U_g2266P608 (.A(G167P74gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2266P608gat) );
AND3XL U_g2272P609 (.A(G164P73gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2272P609gat) );
AND3XL U_g1598P610 (.A(G164P73gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1598P610gat) );
AND3XL U_g1604P611 (.A(G161P72gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1604P611gat) );
AND3XL U_g2278P612 (.A(G161P72gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2278P612gat) );
AND3XL U_g2345P613 (.A(G158P71gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2345P613gat) );
AND3XL U_g1674P614 (.A(G158P71gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1674P614gat) );
AND3XL U_g1680P615 (.A(G152P69gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1680P615gat) );
AND3XL U_g2351P616 (.A(G152P69gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2351P616gat) );
AND3XL U_g2357P617 (.A(G146P67gat), .B(G1691P159gat), .C(G1694P160gat), .Y(G2357P617gat) );
AND3XL U_g1686P618 (.A(G146P67gat), .B(G1689P157gat), .C(G1690P158gat), .Y(G1686P618gat) );
INVXL U_g3724P170_b (.A(G3724P170gat), .Y(G3724P170_bgat) );
AND3XL U_g3734P629 (.A(G123P53gat), .B(G3717P169gat), .C(G3724P170_bgat), .Y(G3734P629gat) );
AND2XL U_g3643P634 (.A(G97P37gat), .B(G4092P176gat), .Y(G3643P634gat) );
AND2XL U_g3637P635 (.A(G97P37gat), .B(G4092P176gat), .Y(G3637P635gat) );
AND2XL U_g3646P636 (.A(G94P36gat), .B(G4092P176gat), .Y(G3646P636gat) );
AND2XL U_g3640P637 (.A(G94P36gat), .B(G4092P176gat), .Y(G3640P637gat) );
INVXL U_g2358P162_b (.A(G2358P162gat), .Y(G2358P162_bgat) );
AND2XL U_g3202P638 (.A(G88P34gat), .B(G2358P162_bgat), .Y(G3202P638gat) );
AND2XL U_g3199P639 (.A(G88P34gat), .B(G2358P162_bgat), .Y(G3199P639gat) );
AND2XL U_g3196P640 (.A(G86P32gat), .B(G2358P162_bgat), .Y(G3196P640gat) );
AND2XL U_g3193P641 (.A(G83P31gat), .B(G2358P162_bgat), .Y(G3193P641gat) );
INVXL U_g210P89_b (.A(G210P89gat), .Y(G210P89_bgat) );
INVXL U_g3548P166_b (.A(G3548P166gat), .Y(G3548P166_bgat) );
AND2XL U_g2592P666 (.A(G210P89_bgat), .B(G3548P166_bgat), .Y(G2592P666gat) );
INVXL U_g218P91_b (.A(G218P91gat), .Y(G218P91_bgat) );
AND2XL U_g2597P667 (.A(G218P91_bgat), .B(G3548P166_bgat), .Y(G2597P667gat) );
INVXL U_g226P93_b (.A(G226P93gat), .Y(G226P93_bgat) );
AND2XL U_g2602P668 (.A(G226P93_bgat), .B(G3548P166_bgat), .Y(G2602P668gat) );
INVXL U_g234P95_b (.A(G234P95gat), .Y(G234P95_bgat) );
AND2XL U_g2607P669 (.A(G234P95_bgat), .B(G3548P166_bgat), .Y(G2607P669gat) );
INVXL U_g257P102_b (.A(G257P102gat), .Y(G257P102_bgat) );
AND2XL U_g2686P670 (.A(G257P102_bgat), .B(G3548P166_bgat), .Y(G2686P670gat) );
INVXL U_g265P104_b (.A(G265P104gat), .Y(G265P104_bgat) );
AND2XL U_g2691P671 (.A(G265P104_bgat), .B(G3548P166_bgat), .Y(G2691P671gat) );
INVXL U_g273P106_b (.A(G273P106gat), .Y(G273P106_bgat) );
AND2XL U_g2696P672 (.A(G273P106_bgat), .B(G3548P166_bgat), .Y(G2696P672gat) );
INVXL U_g281P108_b (.A(G281P108gat), .Y(G281P108_bgat) );
AND2XL U_g2701P673 (.A(G281P108_bgat), .B(G3548P166_bgat), .Y(G2701P673gat) );
INVXL U_g324P120_b (.A(G324P120gat), .Y(G324P120_bgat) );
AND2XL U_g2996P674 (.A(G324P120_bgat), .B(G3548P166_bgat), .Y(G2996P674gat) );
INVXL U_g341P125_b (.A(G341P125gat), .Y(G341P125_bgat) );
AND2XL U_g3003P675 (.A(G341P125_bgat), .B(G3548P166_bgat), .Y(G3003P675gat) );
INVXL U_g351P127_b (.A(G351P127gat), .Y(G351P127_bgat) );
AND2XL U_g3008P676 (.A(G351P127_bgat), .B(G3548P166_bgat), .Y(G3008P676gat) );
AND2XL U_g2869P677 (.A(G2358P162gat), .B(G2822P361_bgat), .Y(G2869P677gat) );
AND2XL U_g2881P678 (.A(G2358P162gat), .B(G2822P361_bgat), .Y(G2881P678gat) );
AND2XL U_g2877P679 (.A(G2358P162gat), .B(G2822P361_bgat), .Y(G2877P679gat) );
AND2XL U_g2873P680 (.A(G2358P162gat), .B(G2822P361_bgat), .Y(G2873P680gat) );
AND2XL U_g2868P681 (.A(G2358P162_bgat), .B(G2822P361_bgat), .Y(G2868P681gat) );
AND2XL U_g2872P682 (.A(G2358P162_bgat), .B(G2822P361_bgat), .Y(G2872P682gat) );
AND2XL U_g2876P683 (.A(G2358P162_bgat), .B(G2822P361_bgat), .Y(G2876P683gat) );
AND2XL U_g2880P684 (.A(G2358P162_bgat), .B(G2822P361_bgat), .Y(G2880P684gat) );
AND3XL U_g3239P685 (.A(G251P100gat), .B(G351P127_bgat), .C(G534P149gat), .Y(G3239P685gat) );
INVXL U_g3550P167_b (.A(G3550P167gat), .Y(G3550P167_bgat) );
AND3XL U_g2990P686 (.A(G351P127_bgat), .B(G534P149gat), .C(G3550P167_bgat), .Y(G2990P686gat) );
AND3XL U_g2984P687 (.A(G341P125_bgat), .B(G523P148gat), .C(G3550P167_bgat), .Y(G2984P687gat) );
AND3XL U_g3235P688 (.A(G251P100gat), .B(G341P125_bgat), .C(G523P148gat), .Y(G3235P688gat) );
AND3XL U_g2975P691 (.A(G324P120_bgat), .B(G503P146gat), .C(G3550P167_bgat), .Y(G2975P691gat) );
AND3XL U_g3229P692 (.A(G251P100gat), .B(G324P120_bgat), .C(G503P146gat), .Y(G3229P692gat) );
INVXL U_g316P118_b (.A(G316P118gat), .Y(G316P118_bgat) );
AND3XL U_g3288P693 (.A(G251P100gat), .B(G316P118_bgat), .C(G490P145gat), .Y(G3288P693gat) );
AND3XL U_g2914P694 (.A(G251P100gat), .B(G316P118_bgat), .C(G490P145gat), .Y(G2914P694gat) );
INVXL U_g308P116_b (.A(G308P116gat), .Y(G308P116_bgat) );
AND3XL U_g2910P695 (.A(G251P100gat), .B(G308P116_bgat), .C(G479P144gat), .Y(G2910P695gat) );
AND3XL U_g3284P696 (.A(G251P100gat), .B(G308P116_bgat), .C(G479P144gat), .Y(G3284P696gat) );
AND3XL U_g3391P697 (.A(G218P91_bgat), .B(G251P100gat), .C(G468P143gat), .Y(G3391P697gat) );
AND3XL U_g2574P698 (.A(G218P91_bgat), .B(G468P143gat), .C(G3550P167_bgat), .Y(G2574P698gat) );
AND3XL U_g3387P699 (.A(G210P89_bgat), .B(G251P100gat), .C(G457P142gat), .Y(G3387P699gat) );
AND3XL U_g2568P700 (.A(G210P89_bgat), .B(G457P142gat), .C(G3550P167_bgat), .Y(G2568P700gat) );
AND3XL U_g3336P701 (.A(G206P87gat), .B(G248P99gat), .C(G446P141gat), .Y(G3336P701gat) );
AND3XL U_g3329P702 (.A(G206P87gat), .B(G248P99gat), .C(G446P141gat), .Y(G3329P702gat) );
AND3XL U_g3399P703 (.A(G234P95_bgat), .B(G251P100gat), .C(G435P140gat), .Y(G3399P703gat) );
AND3XL U_g2586P704 (.A(G234P95_bgat), .B(G435P140gat), .C(G3550P167_bgat), .Y(G2586P704gat) );
AND3XL U_g3395P705 (.A(G226P93_bgat), .B(G251P100gat), .C(G422P139gat), .Y(G3395P705gat) );
AND3XL U_g2580P706 (.A(G226P93_bgat), .B(G422P139gat), .C(G3550P167_bgat), .Y(G2580P706gat) );
AND3XL U_g2674P707 (.A(G273P106_bgat), .B(G411P138gat), .C(G3550P167_bgat), .Y(G2674P707gat) );
AND3XL U_g3065P708 (.A(G251P100gat), .B(G273P106_bgat), .C(G411P138gat), .Y(G3065P708gat) );
AND3XL U_g3061P709 (.A(G251P100gat), .B(G265P104_bgat), .C(G400P137gat), .Y(G3061P709gat) );
AND3XL U_g2668P710 (.A(G265P104_bgat), .B(G400P137gat), .C(G3550P167_bgat), .Y(G2668P710gat) );
AND3XL U_g2662P711 (.A(G257P102_bgat), .B(G389P136gat), .C(G3550P167_bgat), .Y(G2662P711gat) );
AND3XL U_g3057P712 (.A(G251P100gat), .B(G257P102_bgat), .C(G389P136gat), .Y(G3057P712gat) );
AND3XL U_g3069P713 (.A(G251P100gat), .B(G281P108_bgat), .C(G374P134gat), .Y(G3069P713gat) );
AND3XL U_g2680P714 (.A(G281P108_bgat), .B(G374P134gat), .C(G3550P167_bgat), .Y(G2680P714gat) );
INVXL U_g332P122_b (.A(G332P122gat), .Y(G332P122_bgat) );
AND2XL U_g3118P715 (.A(G332P122_bgat), .B(G369P131gat), .Y(G3118P715gat) );
INVXL U_g369P131_b (.A(G369P131gat), .Y(G369P131_bgat) );
OR2XL U_g3422P716 (.A(G361P129gat), .B(G369P131_bgat), .Y(G3422P716gat) );
AND2XL U_g3120P717 (.A(G332P122_bgat), .B(G361P129gat), .Y(G3120P717gat) );
INVXL U_g361P129_b (.A(G361P129gat), .Y(G361P129_bgat) );
OR2XL U_g3423P718 (.A(G361P129_bgat), .B(G369P131gat), .Y(G3423P718gat) );
AND2XL U_g3122P719 (.A(G332P122_bgat), .B(G351P127gat), .Y(G3122P719gat) );
OR2XL U_g3431P720 (.A(G341P125gat), .B(G351P127_bgat), .Y(G3431P720gat) );
AND2XL U_g3124P721 (.A(G332P122_bgat), .B(G341P125gat), .Y(G3124P721gat) );
OR2XL U_g3432P722 (.A(G341P125_bgat), .B(G351P127gat), .Y(G3432P722gat) );
OR2XL U_g3147P723 (.A(G332P122_bgat), .B(G3126P492gat), .Y(G3147P723gat) );
AND2XL U_g3127P724 (.A(G324P120gat), .B(G332P122_bgat), .Y(G3127P724gat) );
AND2XL U_g3129P727 (.A(G316P118gat), .B(G332P122_bgat), .Y(G3129P727gat) );
OR2XL U_g5106P728 (.A(G308P116gat), .B(G316P118_bgat), .Y(G5106P728gat) );
OR2XL U_g5107P729 (.A(G308P116_bgat), .B(G316P118gat), .Y(G5107P729gat) );
AND2XL U_g3131P730 (.A(G308P116gat), .B(G332P122_bgat), .Y(G3131P730gat) );
INVXL U_g302P114_b (.A(G302P114gat), .Y(G302P114_bgat) );
OR2XL U_g5116P731 (.A(G293P112gat), .B(G302P114_bgat), .Y(G5116P731gat) );
AND2XL U_g3133P732 (.A(G302P114gat), .B(G332P122_bgat), .Y(G3133P732gat) );
INVXL U_g293P112_b (.A(G293P112gat), .Y(G293P112_bgat) );
OR2XL U_g5117P735 (.A(G293P112_bgat), .B(G302P114gat), .Y(G5117P735gat) );
AND2XL U_g3135P736 (.A(G293P112gat), .B(G332P122_bgat), .Y(G3135P736gat) );
INVXL U_g335P123_b (.A(G335P123gat), .Y(G335P123_bgat) );
AND2XL U_g2747P737 (.A(G289P110gat), .B(G335P123_bgat), .Y(G2747P737gat) );
INVXL U_g289P110_b (.A(G289P110gat), .Y(G289P110_bgat) );
OR2XL U_g3895P738 (.A(G281P108gat), .B(G289P110_bgat), .Y(G3895P738gat) );
AND2XL U_g2749P739 (.A(G281P108gat), .B(G335P123_bgat), .Y(G2749P739gat) );
OR2XL U_g3896P740 (.A(G281P108_bgat), .B(G289P110gat), .Y(G3896P740gat) );
AND2XL U_g2751P741 (.A(G273P106gat), .B(G335P123_bgat), .Y(G2751P741gat) );
OR2XL U_g3904P742 (.A(G265P104gat), .B(G273P106_bgat), .Y(G3904P742gat) );
AND2XL U_g2753P743 (.A(G265P104gat), .B(G335P123_bgat), .Y(G2753P743gat) );
OR2XL U_g3905P744 (.A(G265P104_bgat), .B(G273P106gat), .Y(G3905P744gat) );
OR2XL U_g3913P745 (.A(G234P95gat), .B(G257P102_bgat), .Y(G3913P745gat) );
AND2XL U_g2755P746 (.A(G257P102gat), .B(G335P123_bgat), .Y(G2755P746gat) );
AND2XL U_g2920P747 (.A(G254P101gat), .B(G293P112_bgat), .Y(G2920P747gat) );
AND2XL U_g2924P748 (.A(G254P101gat), .B(G308P116_bgat), .Y(G2924P748gat) );
AND2XL U_g2929P749 (.A(G254P101gat), .B(G316P118_bgat), .Y(G2929P749gat) );
AND2XL U_g3075P750 (.A(G254P101gat), .B(G257P102_bgat), .Y(G3075P750gat) );
AND2XL U_g3080P751 (.A(G254P101gat), .B(G265P104_bgat), .Y(G3080P751gat) );
AND2XL U_g3085P752 (.A(G254P101gat), .B(G273P106_bgat), .Y(G3085P752gat) );
AND2XL U_g3090P753 (.A(G254P101gat), .B(G281P108_bgat), .Y(G3090P753gat) );
AND2XL U_g3405P754 (.A(G210P89_bgat), .B(G254P101gat), .Y(G3405P754gat) );
AND2XL U_g3410P755 (.A(G218P91_bgat), .B(G254P101gat), .Y(G3410P755gat) );
AND2XL U_g3415P756 (.A(G226P93_bgat), .B(G254P101gat), .Y(G3415P756gat) );
AND2XL U_g3420P757 (.A(G234P95_bgat), .B(G254P101gat), .Y(G3420P757gat) );
AND2XL U_g3244P758 (.A(G254P101gat), .B(G324P120_bgat), .Y(G3244P758gat) );
AND2XL U_g3254P759 (.A(G254P101gat), .B(G351P127_bgat), .Y(G3254P759gat) );
AND2XL U_g3250P760 (.A(G254P101gat), .B(G341P125_bgat), .Y(G3250P760gat) );
AND2XL U_g3293P761 (.A(G254P101gat), .B(G293P112_bgat), .Y(G3293P761gat) );
AND2XL U_g3300P762 (.A(G254P101gat), .B(G316P118_bgat), .Y(G3300P762gat) );
AND2XL U_g3296P763 (.A(G254P101gat), .B(G308P116_bgat), .Y(G3296P763gat) );
AND2XL U_g2907P764 (.A(G251P100gat), .B(G302P114_bgat), .Y(G2907P764gat) );
AND2XL U_g3334P765 (.A(G251P100gat), .B(G361P129_bgat), .Y(G3334P765gat) );
AND2XL U_g3327P766 (.A(G251P100gat), .B(G361P129_bgat), .Y(G3327P766gat) );
AND2XL U_g3281P767 (.A(G251P100gat), .B(G302P114_bgat), .Y(G3281P767gat) );
AND2XL U_g3341P768 (.A(G206P87gat), .B(G242P97gat), .Y(G3341P768gat) );
AND2XL U_g3345P769 (.A(G206P87gat), .B(G242P97gat), .Y(G3345P769gat) );
AND2XL U_g2757P770 (.A(G234P95gat), .B(G335P123_bgat), .Y(G2757P770gat) );
OR2XL U_g3914P771 (.A(G234P95_bgat), .B(G257P102gat), .Y(G3914P771gat) );
OR2XL U_g5364P772 (.A(G218P91gat), .B(G226P93_bgat), .Y(G5364P772gat) );
AND2XL U_g2759P773 (.A(G226P93gat), .B(G335P123_bgat), .Y(G2759P773gat) );
AND2XL U_g2761P774 (.A(G218P91gat), .B(G335P123_bgat), .Y(G2761P774gat) );
OR2XL U_g5365P775 (.A(G218P91_bgat), .B(G226P93gat), .Y(G5365P775gat) );
INVXL U_g206P87_b (.A(G206P87gat), .Y(G206P87_bgat) );
OR2XL U_g5375P776 (.A(G206P87_bgat), .B(G210P89gat), .Y(G5375P776gat) );
AND2XL U_g2763P777 (.A(G210P89gat), .B(G335P123_bgat), .Y(G2763P777gat) );
AND2XL U_g2765P783 (.A(G206P87gat), .B(G335P123_bgat), .Y(G2765P783gat) );
INVXL U_g1691P159_b (.A(G1691P159gat), .Y(G1691P159_bgat) );
AND3XL U_g2259P784 (.A(G203P86gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2259P784gat) );
INVXL U_g1689P157_b (.A(G1689P157gat), .Y(G1689P157_bgat) );
AND3XL U_g1585P785 (.A(G203P86gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1585P785gat) );
AND3XL U_g2253P786 (.A(G200P85gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2253P786gat) );
AND3XL U_g1579P787 (.A(G200P85gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1579P787gat) );
AND3XL U_g2265P788 (.A(G197P84gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2265P788gat) );
AND3XL U_g1591P789 (.A(G197P84gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1591P789gat) );
AND3XL U_g2271P790 (.A(G194P83gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2271P790gat) );
AND3XL U_g1597P791 (.A(G194P83gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1597P791gat) );
AND3XL U_g2277P792 (.A(G191P82gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2277P792gat) );
AND3XL U_g1603P793 (.A(G191P82gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1603P793gat) );
AND3XL U_g1673P794 (.A(G188P81gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1673P794gat) );
AND3XL U_g2344P795 (.A(G188P81gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2344P795gat) );
AND3XL U_g2338P796 (.A(G182P79gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2338P796gat) );
AND3XL U_g1667P797 (.A(G182P79gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1667P797gat) );
AND3XL U_g2331P798 (.A(G176P77gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2331P798gat) );
AND3XL U_g1660P799 (.A(G176P77gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1660P799gat) );
AND3XL U_g2350P800 (.A(G155P70gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2350P800gat) );
AND3XL U_g1679P801 (.A(G155P70gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1679P801gat) );
AND3XL U_g1685P802 (.A(G149P68gat), .B(G1689P157_bgat), .C(G1690P158gat), .Y(G1685P802gat) );
AND3XL U_g2356P803 (.A(G149P68gat), .B(G1691P159_bgat), .C(G1694P160gat), .Y(G2356P803gat) );
AND3XL U_g3838P804 (.A(G131P59gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3838P804gat) );
AND3XL U_g3847P805 (.A(G130P58gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3847P805gat) );
AND3XL U_g3841P806 (.A(G129P57gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3841P806gat) );
AND3XL U_g3789P807 (.A(G128P56gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3789P807gat) );
AND3XL U_g3786P808 (.A(G127P55gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3786P808gat) );
AND3XL U_g3783P809 (.A(G126P54gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3783P809gat) );
AND3XL U_g4081P810 (.A(G123P53gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4081P810gat) );
AND3XL U_g4011P811 (.A(G122P52gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4011P811gat) );
AND3XL U_g4078P812 (.A(G121P51gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4078P812gat) );
AND3XL U_g3844P814 (.A(G119P49gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3844P814gat) );
AND3XL U_g3780P816 (.A(G117P47gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G3780P816gat) );
AND3XL U_g4075P817 (.A(G116P46gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4075P817gat) );
AND3XL U_g4023P818 (.A(G115P45gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4023P818gat) );
AND3XL U_g4020P819 (.A(G114P44gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4020P819gat) );
AND3XL U_g4014P820 (.A(G113P43gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4014P820gat) );
AND3XL U_g4072P821 (.A(G112P42gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4072P821gat) );
AND2XL U_g3195P828 (.A(G87P33gat), .B(G2358P162gat), .Y(G3195P828gat) );
AND2XL U_g3192P829 (.A(G83P31gat), .B(G2358P162gat), .Y(G3192P829gat) );
AND3XL U_g4017P836 (.A(G53P19gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4017P836gat) );
AND3XL U_g4069P837 (.A(G52P18gat), .B(G4091P175_bgat), .C(G4092P176gat), .Y(G4069P837gat) );
AND2XL U_g3201P842 (.A(G34P12gat), .B(G2358P162gat), .Y(G3201P842gat) );
AND2XL U_g3198P843 (.A(G34P12gat), .B(G2358P162gat), .Y(G3198P843gat) );
OR3XL U_g3255P854 (.A(G534P149gat), .B(G3253P480gat), .C(G3254P759gat), .Y(G3255P854gat) );
OR2XL U_g3240P855 (.A(G3238P409gat), .B(G3239P685gat), .Y(G3240P855gat) );
OR3XL U_g3009P856 (.A(G534P149gat), .B(G3006P396gat), .C(G3008P676gat), .Y(G3009P856gat) );
OR2XL U_g2991P857 (.A(G2988P410gat), .B(G2990P686gat), .Y(G2991P857gat) );
OR2XL U_g2985P858 (.A(G2982P413gat), .B(G2984P687gat), .Y(G2985P858gat) );
OR3XL U_g3004P859 (.A(G523P148gat), .B(G3001P395gat), .C(G3003P675gat), .Y(G3004P859gat) );
OR2XL U_g3236P860 (.A(G3234P414gat), .B(G3235P688gat), .Y(G3236P860gat) );
OR3XL U_g3251P861 (.A(G523P148gat), .B(G3249P486gat), .C(G3250P760gat), .Y(G3251P861gat) );
INVXL U_g3232P418_b (.A(G3232P418gat), .Y(G3232P418_bgat) );
AND2XL U_g5307P862 (.A(G3247P417gat), .B(G3232P418_bgat), .Y(G5307P862gat) );
INVXL U_g2979P420_b (.A(G2979P420gat), .Y(G2979P420_bgat) );
AND2XL U_g3015P863 (.A(G2999P419gat), .B(G2979P420_bgat), .Y(G3015P863gat) );
AND2XL U_g2036P864 (.A(G514P147gat), .B(G3147P723gat), .Y(G2036P864gat) );
AND2XL U_g1789P865 (.A(G514P147gat), .B(G3147P723gat), .Y(G1789P865gat) );
OR2XL U_g2976P866 (.A(G2973P423gat), .B(G2975P691gat), .Y(G2976P866gat) );
OR3XL U_g2997P867 (.A(G503P146gat), .B(G2994P394gat), .C(G2996P674gat), .Y(G2997P867gat) );
OR2XL U_g3230P868 (.A(G3228P424gat), .B(G3229P692gat), .Y(G3230P868gat) );
OR3XL U_g3245P869 (.A(G503P146gat), .B(G3243P498gat), .C(G3244P758gat), .Y(G3245P869gat) );
OR3XL U_g3301P870 (.A(G490P145gat), .B(G3299P507gat), .C(G3300P762gat), .Y(G3301P870gat) );
OR2XL U_g3289P871 (.A(G3287P427gat), .B(G3288P693gat), .Y(G3289P871gat) );
OR3XL U_g2930P872 (.A(G490P145gat), .B(G2927P510gat), .C(G2929P749gat), .Y(G2930P872gat) );
OR2XL U_g2915P873 (.A(G2913P428gat), .B(G2914P694gat), .Y(G2915P873gat) );
OR2XL U_g2911P874 (.A(G2909P431gat), .B(G2910P695gat), .Y(G2911P874gat) );
OR3XL U_g2925P875 (.A(G479P144gat), .B(G2922P518gat), .C(G2924P748gat), .Y(G2925P875gat) );
OR2XL U_g3285P876 (.A(G3283P432gat), .B(G3284P696gat), .Y(G3285P876gat) );
OR3XL U_g3297P877 (.A(G479P144gat), .B(G3295P515gat), .C(G3296P763gat), .Y(G3297P877gat) );
OR3XL U_g3411P878 (.A(G468P143gat), .B(G3408P566gat), .C(G3410P755gat), .Y(G3411P878gat) );
OR2XL U_g3392P879 (.A(G3390P435gat), .B(G3391P697gat), .Y(G3392P879gat) );
OR3XL U_g2598P880 (.A(G468P143gat), .B(G2595P387gat), .C(G2597P667gat), .Y(G2598P880gat) );
OR2XL U_g2575P881 (.A(G2572P436gat), .B(G2574P698gat), .Y(G2575P881gat) );
OR2XL U_g3388P882 (.A(G3386P439gat), .B(G3387P699gat), .Y(G3388P882gat) );
OR3XL U_g3406P883 (.A(G457P142gat), .B(G3403P565gat), .C(G3405P754gat), .Y(G3406P883gat) );
OR2XL U_g2569P884 (.A(G2566P440gat), .B(G2568P700gat), .Y(G2569P884gat) );
OR3XL U_g2593P885 (.A(G457P142gat), .B(G2590P386gat), .C(G2592P666gat), .Y(G2593P885gat) );
AND3XL U_g3337P886 (.A(G206P87_bgat), .B(G251P100gat), .C(G446P141gat), .Y(G3337P886gat) );
AND3XL U_g3330P887 (.A(G206P87_bgat), .B(G251P100gat), .C(G446P141gat), .Y(G3330P887gat) );
OR3XL U_g3421P888 (.A(G435P140gat), .B(G3418P568gat), .C(G3420P757gat), .Y(G3421P888gat) );
OR2XL U_g3400P889 (.A(G3398P445gat), .B(G3399P703gat), .Y(G3400P889gat) );
OR3XL U_g2608P890 (.A(G435P140gat), .B(G2605P389gat), .C(G2607P669gat), .Y(G2608P890gat) );
OR2XL U_g2587P891 (.A(G2584P446gat), .B(G2586P704gat), .Y(G2587P891gat) );
OR2XL U_g3396P892 (.A(G3394P449gat), .B(G3395P705gat), .Y(G3396P892gat) );
OR3XL U_g3416P893 (.A(G422P139gat), .B(G3413P567gat), .C(G3415P756gat), .Y(G3416P893gat) );
OR2XL U_g2581P894 (.A(G2578P450gat), .B(G2580P706gat), .Y(G2581P894gat) );
OR3XL U_g2603P895 (.A(G422P139gat), .B(G2600P388gat), .C(G2602P668gat), .Y(G2603P895gat) );
OR2XL U_g2675P896 (.A(G2672P453gat), .B(G2674P707gat), .Y(G2675P896gat) );
OR3XL U_g2697P897 (.A(G411P138gat), .B(G2694P392gat), .C(G2696P672gat), .Y(G2697P897gat) );
OR2XL U_g3066P898 (.A(G3064P454gat), .B(G3065P708gat), .Y(G3066P898gat) );
OR3XL U_g3086P899 (.A(G411P138gat), .B(G3083P545gat), .C(G3085P752gat), .Y(G3086P899gat) );
OR3XL U_g3081P900 (.A(G400P137gat), .B(G3078P553gat), .C(G3080P751gat), .Y(G3081P900gat) );
OR2XL U_g3062P901 (.A(G3060P457gat), .B(G3061P709gat), .Y(G3062P901gat) );
OR3XL U_g2692P902 (.A(G400P137gat), .B(G2689P391gat), .C(G2691P671gat), .Y(G2692P902gat) );
OR2XL U_g2669P903 (.A(G2666P458gat), .B(G2668P710gat), .Y(G2669P903gat) );
OR2XL U_g2663P904 (.A(G2660P461gat), .B(G2662P711gat), .Y(G2663P904gat) );
OR3XL U_g2687P905 (.A(G389P136gat), .B(G2684P390gat), .C(G2686P670gat), .Y(G2687P905gat) );
OR2XL U_g3058P906 (.A(G3056P462gat), .B(G3057P712gat), .Y(G3058P906gat) );
OR3XL U_g3076P907 (.A(G389P136gat), .B(G3073P560gat), .C(G3075P750gat), .Y(G3076P907gat) );
OR3XL U_g3091P908 (.A(G374P134gat), .B(G3088P539gat), .C(G3090P753gat), .Y(G3091P908gat) );
OR2XL U_g3070P909 (.A(G3068P466gat), .B(G3069P713gat), .Y(G3070P909gat) );
OR3XL U_g2702P910 (.A(G374P134gat), .B(G2699P393gat), .C(G2701P673gat), .Y(G2702P910gat) );
OR2XL U_g2681P911 (.A(G2678P467gat), .B(G2680P714gat), .Y(G2681P911gat) );
OR2XL U_g5126P912 (.A(G3119P470gat), .B(G3118P715gat), .Y(G5126P912gat) );
INVXL U_g3422P716_b (.A(G3422P716gat), .Y(G3422P716_bgat) );
INVXL U_g3423P718_b (.A(G3423P718gat), .Y(G3423P718_bgat) );
OR2XL U_g3424P913 (.A(G3422P716_bgat), .B(G3423P718_bgat), .Y(G3424P913gat) );
OR2XL U_g3137P914 (.A(G3121P472gat), .B(G3120P717gat), .Y(G3137P914gat) );
OR2XL U_g3335P915 (.A(G3333P473gat), .B(G3334P765gat), .Y(G3335P915gat) );
OR2XL U_g3328P916 (.A(G3326P475gat), .B(G3327P766gat), .Y(G3328P916gat) );
OR2XL U_g3139P917 (.A(G3123P478gat), .B(G3122P719gat), .Y(G3139P917gat) );
INVXL U_g3431P720_b (.A(G3431P720gat), .Y(G3431P720_bgat) );
INVXL U_g3432P722_b (.A(G3432P722gat), .Y(G3432P722_bgat) );
OR2XL U_g3433P918 (.A(G3431P720_bgat), .B(G3432P722_bgat), .Y(G3433P918gat) );
OR2XL U_g3143P919 (.A(G3125P485gat), .B(G3124P721gat), .Y(G3143P919gat) );
OR2XL U_g3151P923 (.A(G3128P497gat), .B(G3127P724gat), .Y(G3151P923gat) );
OR2XL U_g3155P924 (.A(G3130P505gat), .B(G3129P727gat), .Y(G3155P924gat) );
INVXL U_g5106P728_b (.A(G5106P728gat), .Y(G5106P728_bgat) );
INVXL U_g5107P729_b (.A(G5107P729gat), .Y(G5107P729_bgat) );
OR2XL U_g5209P925 (.A(G5106P728_bgat), .B(G5107P729_bgat), .Y(G5209P925gat) );
OR2XL U_g3161P926 (.A(G3132P513gat), .B(G3131P730gat), .Y(G3161P926gat) );
OR2XL U_g3165P927 (.A(G3134P521gat), .B(G3133P732gat), .Y(G3165P927gat) );
OR2XL U_g3282P928 (.A(G3280P522gat), .B(G3281P767gat), .Y(G3282P928gat) );
INVXL U_g5116P731_b (.A(G5116P731gat), .Y(G5116P731_bgat) );
INVXL U_g5117P735_b (.A(G5117P735gat), .Y(G5117P735_bgat) );
OR2XL U_g5206P929 (.A(G5116P731_bgat), .B(G5117P735_bgat), .Y(G5206P929gat) );
OR2XL U_g2908P930 (.A(G2906P525gat), .B(G2907P764gat), .Y(G2908P930gat) );
OR2XL U_g3167P931 (.A(G3136P529gat), .B(G3135P736gat), .Y(G3167P931gat) );
OR2XL U_g5322P932 (.A(G3292P531gat), .B(G3293P761gat), .Y(G5322P932gat) );
OR2XL U_g2933P933 (.A(G2918P533gat), .B(G2920P747gat), .Y(G2933P933gat) );
OR2XL U_g5178P934 (.A(G2748P535gat), .B(G2747P737gat), .Y(G5178P934gat) );
INVXL U_g3895P738_b (.A(G3895P738gat), .Y(G3895P738_bgat) );
INVXL U_g3896P740_b (.A(G3896P740gat), .Y(G3896P740_bgat) );
OR2XL U_g3897P935 (.A(G3895P738_bgat), .B(G3896P740_bgat), .Y(G3897P935gat) );
OR2XL U_g2767P936 (.A(G2750P537gat), .B(G2749P739gat), .Y(G2767P936gat) );
OR2XL U_g2772P937 (.A(G2752P544gat), .B(G2751P741gat), .Y(G2772P937gat) );
INVXL U_g3904P742_b (.A(G3904P742gat), .Y(G3904P742_bgat) );
INVXL U_g3905P744_b (.A(G3905P744gat), .Y(G3905P744_bgat) );
OR2XL U_g3906P938 (.A(G3904P742_bgat), .B(G3905P744_bgat), .Y(G3906P938gat) );
OR2XL U_g2776P939 (.A(G2754P551gat), .B(G2753P743gat), .Y(G2776P939gat) );
OR2XL U_g2780P940 (.A(G2756P558gat), .B(G2755P746gat), .Y(G2780P940gat) );
INVXL U_g3913P745_b (.A(G3913P745gat), .Y(G3913P745_bgat) );
INVXL U_g3914P771_b (.A(G3914P771gat), .Y(G3914P771_bgat) );
OR2XL U_g3915P941 (.A(G3913P745_bgat), .B(G3914P771_bgat), .Y(G3915P941gat) );
AND2XL U_g3342P942 (.A(G206P87_bgat), .B(G254P101gat), .Y(G3342P942gat) );
AND2XL U_g3346P943 (.A(G206P87_bgat), .B(G254P101gat), .Y(G3346P943gat) );
OR2XL U_g2784P944 (.A(G2758P569gat), .B(G2757P770gat), .Y(G2784P944gat) );
OR2XL U_g2788P945 (.A(G2760P575gat), .B(G2759P773gat), .Y(G2788P945gat) );
INVXL U_g5364P772_b (.A(G5364P772gat), .Y(G5364P772_bgat) );
INVXL U_g5365P775_b (.A(G5365P775gat), .Y(G5365P775_bgat) );
OR2XL U_g5399P946 (.A(G5364P772_bgat), .B(G5365P775_bgat), .Y(G5399P946gat) );
OR2XL U_g2794P947 (.A(G2762P581gat), .B(G2761P774gat), .Y(G2794P947gat) );
OR2XL U_g2798P948 (.A(G2764P587gat), .B(G2763P777gat), .Y(G2798P948gat) );
OR2XL U_g5374P949 (.A(G206P87gat), .B(G210P89_bgat), .Y(G5374P949gat) );
OR2XL U_g2802P950 (.A(G2766P593gat), .B(G2765P783gat), .Y(G2802P950gat) );
OR2XL U_g3203P951 (.A(G3202P638gat), .B(G3201P842gat), .Y(G3203P951gat) );
OR2XL U_g3200P952 (.A(G3199P639gat), .B(G3198P843gat), .Y(G3200P952gat) );
OR2XL U_g3197P953 (.A(G3196P640gat), .B(G3195P828gat), .Y(G3197P953gat) );
OR2XL U_g3194P954 (.A(G3193P641gat), .B(G3192P829gat), .Y(G3194P954gat) );
AND3XL U_g2870P955 (.A(G82P30gat), .B(G2358P162_bgat), .C(G2822P361gat), .Y(G2870P955gat) );
AND3XL U_g2875P956 (.A(G81P29gat), .B(G2358P162gat), .C(G2822P361gat), .Y(G2875P956gat) );
AND3XL U_g2871P957 (.A(G80P28gat), .B(G2358P162gat), .C(G2822P361gat), .Y(G2871P957gat) );
AND3XL U_g2866P958 (.A(G79P27gat), .B(G2358P162_bgat), .C(G2822P361gat), .Y(G2866P958gat) );
AND3XL U_g2874P959 (.A(G26P9gat), .B(G2358P162_bgat), .C(G2822P361gat), .Y(G2874P959gat) );
AND3XL U_g2879P960 (.A(G25P8gat), .B(G2358P162gat), .C(G2822P361gat), .Y(G2879P960gat) );
AND3XL U_g2878P961 (.A(G24P7gat), .B(G2358P162_bgat), .C(G2822P361gat), .Y(G2878P961gat) );
AND3XL U_g2867P962 (.A(G23P6gat), .B(G2358P162gat), .C(G2822P361gat), .Y(G2867P962gat) );
AND3XL U_g3845P963 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3015P863gat), .Y(G3845P963gat) );
AND2XL U_g2081P970 (.A(G534P149gat), .B(G3139P917gat), .Y(G2081P970gat) );
AND2XL U_g1823P971 (.A(G534P149gat), .B(G3139P917gat), .Y(G1823P971gat) );
AND2XL U_g1806P974 (.A(G523P148gat), .B(G3143P919gat), .Y(G1806P974gat) );
AND2XL U_g2059P975 (.A(G523P148gat), .B(G3143P919gat), .Y(G2059P975gat) );
INVXL U_g3147P723_b (.A(G3147P723gat), .Y(G3147P723_bgat) );
OR2XL U_g2019P978 (.A(G514P147gat), .B(G3147P723_bgat), .Y(G2019P978gat) );
OR2XL U_g1777P979 (.A(G514P147gat), .B(G3147P723_bgat), .Y(G1777P979gat) );
AND2XL U_g2018P982 (.A(G503P146gat), .B(G3151P923gat), .Y(G2018P982gat) );
AND2XL U_g1775P983 (.A(G503P146gat), .B(G3151P923gat), .Y(G1775P983gat) );
INVXL U_g490P145_b (.A(G490P145gat), .Y(G490P145_bgat) );
INVXL U_g3155P924_b (.A(G3155P924gat), .Y(G3155P924_bgat) );
AND2XL U_g4812P986 (.A(G490P145_bgat), .B(G3155P924_bgat), .Y(G4812P986gat) );
AND2XL U_g2001P987 (.A(G490P145gat), .B(G3155P924gat), .Y(G2001P987gat) );
AND2XL U_g1749P988 (.A(G490P145gat), .B(G3155P924gat), .Y(G1749P988gat) );
AND2XL U_g4716P989 (.A(G490P145_bgat), .B(G3155P924_bgat), .Y(G4716P989gat) );
AND2XL U_g1742P992 (.A(G479P144gat), .B(G3161P926gat), .Y(G1742P992gat) );
AND2XL U_g1995P993 (.A(G479P144gat), .B(G3161P926gat), .Y(G1995P993gat) );
AND2XL U_g1064P996 (.A(G468P143gat), .B(G2794P947gat), .Y(G1064P996gat) );
AND2XL U_g1318P997 (.A(G468P143gat), .B(G2794P947gat), .Y(G1318P997gat) );
AND2XL U_g1301P1000 (.A(G457P142gat), .B(G2798P948gat), .Y(G1301P1000gat) );
AND2XL U_g1046P1001 (.A(G457P142gat), .B(G2798P948gat), .Y(G1046P1001gat) );
OR3XL U_g3347P1002 (.A(G446P141gat), .B(G3345P769gat), .C(G3346P943gat), .Y(G3347P1002gat) );
OR2XL U_g3338P1003 (.A(G3336P701gat), .B(G3337P886gat), .Y(G3338P1003gat) );
OR3XL U_g3343P1004 (.A(G446P141gat), .B(G3341P768gat), .C(G3342P942gat), .Y(G3343P1004gat) );
OR2XL U_g3331P1005 (.A(G3329P702gat), .B(G3330P887gat), .Y(G3331P1005gat) );
AND2XL U_g1031P1006 (.A(G446P141gat), .B(G2802P950gat), .Y(G1031P1006gat) );
AND2XL U_g1286P1007 (.A(G446P141gat), .B(G2802P950gat), .Y(G1286P1007gat) );
AND2XL U_g1341P1010 (.A(G435P140gat), .B(G2784P944gat), .Y(G1341P1010gat) );
AND2XL U_g1097P1011 (.A(G435P140gat), .B(G2784P944gat), .Y(G1097P1011gat) );
AND2XL U_g1071P1014 (.A(G422P139gat), .B(G2788P945gat), .Y(G1071P1014gat) );
INVXL U_g422P139_b (.A(G422P139gat), .Y(G422P139_bgat) );
INVXL U_g2788P945_b (.A(G2788P945gat), .Y(G2788P945_bgat) );
AND2XL U_g4228P1015 (.A(G422P139_bgat), .B(G2788P945_bgat), .Y(G4228P1015gat) );
AND2XL U_g4348P1016 (.A(G422P139_bgat), .B(G2788P945_bgat), .Y(G4348P1016gat) );
AND2XL U_g1324P1017 (.A(G422P139gat), .B(G2788P945gat), .Y(G1324P1017gat) );
AND2XL U_g1145P1020 (.A(G411P138gat), .B(G2772P937gat), .Y(G1145P1020gat) );
AND2XL U_g1404P1021 (.A(G411P138gat), .B(G2772P937gat), .Y(G1404P1021gat) );
AND2XL U_g1382P1024 (.A(G400P137gat), .B(G2776P939gat), .Y(G1382P1024gat) );
AND2XL U_g1128P1025 (.A(G400P137gat), .B(G2776P939gat), .Y(G1128P1025gat) );
AND2XL U_g1111P1028 (.A(G389P136gat), .B(G2780P940gat), .Y(G1111P1028gat) );
AND2XL U_g1359P1029 (.A(G389P136gat), .B(G2780P940gat), .Y(G1359P1029gat) );
INVXL U_g374P134_b (.A(G374P134gat), .Y(G374P134_bgat) );
INVXL U_g2767P936_b (.A(G2767P936gat), .Y(G2767P936_bgat) );
AND2XL U_g4464P1032 (.A(G374P134_bgat), .B(G2767P936_bgat), .Y(G4464P1032gat) );
AND2XL U_g1412P1033 (.A(G374P134gat), .B(G2767P936gat), .Y(G1412P1033gat) );
AND2XL U_g1160P1034 (.A(G374P134gat), .B(G2767P936gat), .Y(G1160P1034gat) );
AND3XL U_g3514P1057 (.A(G324P120_bgat), .B(G3424P913gat), .C(G3433P918gat), .Y(G3514P1057gat) );
INVXL U_g5375P776_b (.A(G5375P776gat), .Y(G5375P776_bgat) );
INVXL U_g5374P949_b (.A(G5374P949gat), .Y(G5374P949_bgat) );
OR2XL U_g5396P1110 (.A(G5375P776_bgat), .B(G5374P949_bgat), .Y(G5396P1110gat) );
INVXL U_g2908P930_b (.A(G2908P930gat), .Y(G2908P930_bgat) );
AND3XL U_g4076P1118 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2908P930_bgat), .Y(G4076P1118gat) );
AND3XL U_g4079P1119 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2933P933gat), .Y(G4079P1119gat) );
INVXL U_g3335P915_b (.A(G3335P915gat), .Y(G3335P915_bgat) );
AND3XL U_g3836P1120 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3335P915_bgat), .Y(G3836P1120gat) );
INVXL U_g3717P169_b (.A(G3717P169gat), .Y(G3717P169_bgat) );
AND3XL U_g3731P1121 (.A(G3717P169_bgat), .B(G3724P170_bgat), .C(G2933P933gat), .Y(G3731P1121gat) );
INVXL U_g3240P855_b (.A(G3240P855gat), .Y(G3240P855_bgat) );
AND2XL U_g5299P1122 (.A(G3255P854gat), .B(G3240P855_bgat), .Y(G5299P1122gat) );
INVXL U_g2991P857_b (.A(G2991P857gat), .Y(G2991P857_bgat) );
AND2XL U_g3021P1123 (.A(G3009P856gat), .B(G2991P857_bgat), .Y(G3021P1123gat) );
INVXL U_g3139P917_b (.A(G3139P917gat), .Y(G3139P917_bgat) );
OR2XL U_g2065P1124 (.A(G534P149gat), .B(G3139P917_bgat), .Y(G2065P1124gat) );
OR2XL U_g1811P1125 (.A(G534P149gat), .B(G3139P917_bgat), .Y(G1811P1125gat) );
INVXL U_g2985P858_b (.A(G2985P858gat), .Y(G2985P858_bgat) );
AND2XL U_g3018P1126 (.A(G2985P858_bgat), .B(G3004P859gat), .Y(G3018P1126gat) );
INVXL U_g3236P860_b (.A(G3236P860gat), .Y(G3236P860_bgat) );
AND2XL U_g5296P1127 (.A(G3236P860_bgat), .B(G3251P861gat), .Y(G5296P1127gat) );
INVXL U_g3143P919_b (.A(G3143P919gat), .Y(G3143P919_bgat) );
OR2XL U_g1793P1128 (.A(G523P148gat), .B(G3143P919_bgat), .Y(G1793P1128gat) );
OR2XL U_g2040P1129 (.A(G523P148gat), .B(G3143P919_bgat), .Y(G2040P1129gat) );
INVXL U_g514P147_b (.A(G514P147gat), .Y(G514P147_bgat) );
OR2XL U_g2020P1130 (.A(G514P147_bgat), .B(G3147P723gat), .Y(G2020P1130gat) );
OR2XL U_g1776P1131 (.A(G514P147_bgat), .B(G3147P723gat), .Y(G1776P1131gat) );
INVXL U_g2976P866_b (.A(G2976P866gat), .Y(G2976P866_bgat) );
AND2XL U_g3012P1132 (.A(G2976P866_bgat), .B(G2997P867gat), .Y(G3012P1132gat) );
INVXL U_g3230P868_b (.A(G3230P868gat), .Y(G3230P868_bgat) );
AND2XL U_g5304P1133 (.A(G3230P868_bgat), .B(G3245P869gat), .Y(G5304P1133gat) );
INVXL U_g3151P923_b (.A(G3151P923gat), .Y(G3151P923_bgat) );
OR2XL U_g2007P1134 (.A(G503P146gat), .B(G3151P923_bgat), .Y(G2007P1134gat) );
OR2XL U_g1766P1135 (.A(G503P146gat), .B(G3151P923_bgat), .Y(G1766P1135gat) );
INVXL U_g3289P871_b (.A(G3289P871gat), .Y(G3289P871_bgat) );
AND2XL U_g5315P1136 (.A(G3301P870gat), .B(G3289P871_bgat), .Y(G5315P1136gat) );
INVXL U_g2915P873_b (.A(G2915P873gat), .Y(G2915P873_bgat) );
AND2XL U_g2942P1137 (.A(G2930P872gat), .B(G2915P873_bgat), .Y(G2942P1137gat) );
OR2XL U_g2097P1138 (.A(G490P145gat), .B(G3155P924_bgat), .Y(G2097P1138gat) );
OR2XL U_g1757P1141 (.A(G490P145gat), .B(G3155P924_bgat), .Y(G1757P1141gat) );
INVXL U_g2911P874_b (.A(G2911P874gat), .Y(G2911P874_bgat) );
AND2XL U_g2939P1144 (.A(G2911P874_bgat), .B(G2925P875gat), .Y(G2939P1144gat) );
INVXL U_g3285P876_b (.A(G3285P876gat), .Y(G3285P876_bgat) );
AND2XL U_g5312P1145 (.A(G3285P876_bgat), .B(G3297P877gat), .Y(G5312P1145gat) );
INVXL U_g3161P926_b (.A(G3161P926gat), .Y(G3161P926_bgat) );
OR2XL U_g1729P1146 (.A(G479P144gat), .B(G3161P926_bgat), .Y(G1729P1146gat) );
AND3XL U_g1846P1147 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G1742P992gat), .Y(G1846P1147gat) );
AND2XL U_g1849P1148 (.A(G3165P927_bgat), .B(G1742P992gat), .Y(G1849P1148gat) );
AND2XL U_g1852P1149 (.A(G3165P927_bgat), .B(G1742P992gat), .Y(G1852P1149gat) );
OR2XL U_g1982P1150 (.A(G479P144gat), .B(G3161P926_bgat), .Y(G1982P1150gat) );
AND2XL U_g2122P1151 (.A(G3165P927_bgat), .B(G1995P993gat), .Y(G2122P1151gat) );
AND3XL U_g2116P1152 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G1995P993gat), .Y(G2116P1152gat) );
AND2XL U_g2119P1153 (.A(G3165P927_bgat), .B(G1995P993gat), .Y(G2119P1153gat) );
INVXL U_g3392P879_b (.A(G3392P879gat), .Y(G3392P879_bgat) );
AND2XL U_g5276P1154 (.A(G3411P878gat), .B(G3392P879_bgat), .Y(G5276P1154gat) );
INVXL U_g2575P881_b (.A(G2575P881gat), .Y(G2575P881_bgat) );
AND2XL U_g2615P1155 (.A(G2598P880gat), .B(G2575P881_bgat), .Y(G2615P1155gat) );
INVXL U_g2794P947_b (.A(G2794P947gat), .Y(G2794P947_bgat) );
OR2XL U_g1051P1156 (.A(G468P143gat), .B(G2794P947_bgat), .Y(G1051P1156gat) );
OR2XL U_g1305P1157 (.A(G468P143gat), .B(G2794P947_bgat), .Y(G1305P1157gat) );
INVXL U_g3388P882_b (.A(G3388P882gat), .Y(G3388P882_bgat) );
AND2XL U_g5289P1158 (.A(G3388P882_bgat), .B(G3406P883gat), .Y(G5289P1158gat) );
INVXL U_g2569P884_b (.A(G2569P884gat), .Y(G2569P884_bgat) );
AND2XL U_g2611P1159 (.A(G2569P884_bgat), .B(G2593P885gat), .Y(G2611P1159gat) );
INVXL U_g2798P948_b (.A(G2798P948gat), .Y(G2798P948_bgat) );
OR2XL U_g1287P1160 (.A(G457P142gat), .B(G2798P948_bgat), .Y(G1287P1160gat) );
OR2XL U_g1033P1161 (.A(G457P142gat), .B(G2798P948_bgat), .Y(G1033P1161gat) );
INVXL U_g2802P950_b (.A(G2802P950gat), .Y(G2802P950_bgat) );
OR2XL U_g1022P1164 (.A(G446P141gat), .B(G2802P950_bgat), .Y(G1022P1164gat) );
OR2XL U_g1276P1165 (.A(G446P141gat), .B(G2802P950_bgat), .Y(G1276P1165gat) );
INVXL U_g3400P889_b (.A(G3400P889gat), .Y(G3400P889_bgat) );
AND2XL U_g5268P1166 (.A(G3421P888gat), .B(G3400P889_bgat), .Y(G5268P1166gat) );
INVXL U_g2587P891_b (.A(G2587P891gat), .Y(G2587P891_bgat) );
AND2XL U_g2623P1167 (.A(G2608P890gat), .B(G2587P891_bgat), .Y(G2623P1167gat) );
INVXL U_g2784P944_b (.A(G2784P944gat), .Y(G2784P944_bgat) );
OR2XL U_g1330P1168 (.A(G435P140gat), .B(G2784P944_bgat), .Y(G1330P1168gat) );
OR2XL U_g1088P1169 (.A(G435P140gat), .B(G2784P944_bgat), .Y(G1088P1169gat) );
INVXL U_g3396P892_b (.A(G3396P892gat), .Y(G3396P892_bgat) );
AND2XL U_g5279P1170 (.A(G3396P892_bgat), .B(G3416P893gat), .Y(G5279P1170gat) );
INVXL U_g2581P894_b (.A(G2581P894gat), .Y(G2581P894_bgat) );
AND2XL U_g2619P1171 (.A(G2581P894_bgat), .B(G2603P895gat), .Y(G2619P1171gat) );
OR2XL U_g1079P1172 (.A(G422P139gat), .B(G2788P945_bgat), .Y(G1079P1172gat) );
OR2XL U_g1420P1175 (.A(G422P139gat), .B(G2788P945_bgat), .Y(G1420P1175gat) );
INVXL U_g2675P896_b (.A(G2675P896gat), .Y(G2675P896_bgat) );
AND2XL U_g2713P1178 (.A(G2675P896_bgat), .B(G2697P897gat), .Y(G2713P1178gat) );
INVXL U_g3066P898_b (.A(G3066P898gat), .Y(G3066P898_bgat) );
AND2XL U_g5263P1179 (.A(G3066P898_bgat), .B(G3086P899gat), .Y(G5263P1179gat) );
INVXL U_g2772P937_b (.A(G2772P937gat), .Y(G2772P937_bgat) );
OR2XL U_g1133P1180 (.A(G411P138gat), .B(G2772P937_bgat), .Y(G1133P1180gat) );
OR2XL U_g1388P1181 (.A(G411P138gat), .B(G2772P937_bgat), .Y(G1388P1181gat) );
INVXL U_g3062P901_b (.A(G3062P901gat), .Y(G3062P901_bgat) );
AND2XL U_g5260P1182 (.A(G3081P900gat), .B(G3062P901_bgat), .Y(G5260P1182gat) );
INVXL U_g2669P903_b (.A(G2669P903gat), .Y(G2669P903_bgat) );
AND2XL U_g2709P1183 (.A(G2692P902gat), .B(G2669P903_bgat), .Y(G2709P1183gat) );
INVXL U_g2776P939_b (.A(G2776P939gat), .Y(G2776P939_bgat) );
OR2XL U_g1363P1184 (.A(G400P137gat), .B(G2776P939_bgat), .Y(G1363P1184gat) );
OR2XL U_g1115P1185 (.A(G400P137gat), .B(G2776P939_bgat), .Y(G1115P1185gat) );
INVXL U_g2663P904_b (.A(G2663P904gat), .Y(G2663P904_bgat) );
AND2XL U_g2705P1186 (.A(G2663P904_bgat), .B(G2687P905gat), .Y(G2705P1186gat) );
INVXL U_g3058P906_b (.A(G3058P906gat), .Y(G3058P906_bgat) );
AND2XL U_g5271P1187 (.A(G3058P906_bgat), .B(G3076P907gat), .Y(G5271P1187gat) );
INVXL U_g2780P940_b (.A(G2780P940gat), .Y(G2780P940_bgat) );
OR2XL U_g1099P1188 (.A(G389P136gat), .B(G2780P940_bgat), .Y(G1099P1188gat) );
OR2XL U_g1342P1189 (.A(G389P136gat), .B(G2780P940_bgat), .Y(G1342P1189gat) );
INVXL U_g3070P909_b (.A(G3070P909gat), .Y(G3070P909_bgat) );
AND2XL U_g3852P1190 (.A(G3091P908gat), .B(G3070P909_bgat), .Y(G3852P1190gat) );
INVXL U_g2681P911_b (.A(G2681P911gat), .Y(G2681P911_bgat) );
AND2XL U_g2717P1191 (.A(G2702P910gat), .B(G2681P911_bgat), .Y(G2717P1191gat) );
OR2XL U_g1428P1192 (.A(G374P134gat), .B(G2767P936_bgat), .Y(G1428P1192gat) );
OR2XL U_g1151P1195 (.A(G374P134gat), .B(G2767P936_bgat), .Y(G1151P1195gat) );
OR2XL U_g3452P1196 (.A(G5126P912gat), .B(G3137P914_bgat), .Y(G3452P1196gat) );
OR2XL U_g3462P1210 (.A(G3147P723gat), .B(G3151P923_bgat), .Y(G3462P1210gat) );
INVXL U_g3424P913_b (.A(G3424P913gat), .Y(G3424P913_bgat) );
INVXL U_g3433P918_b (.A(G3433P918gat), .Y(G3433P918_bgat) );
AND3XL U_g3517P1214 (.A(G324P120_bgat), .B(G3424P913_bgat), .C(G3433P918_bgat), .Y(G3517P1214gat) );
AND3XL U_g3516P1215 (.A(G324P120gat), .B(G3424P913gat), .C(G3433P918_bgat), .Y(G3516P1215gat) );
AND3XL U_g3513P1216 (.A(G324P120gat), .B(G3424P913_bgat), .C(G3433P918gat), .Y(G3513P1216gat) );
INVXL U_g5209P925_b (.A(G5209P925gat), .Y(G5209P925_bgat) );
OR2XL U_g5214P1220 (.A(G5209P925_bgat), .B(G5206P929gat), .Y(G5214P1220gat) );
AND2XL U_g1845P1226 (.A(G3165P927gat), .B(G3167P931_bgat), .Y(G1845P1226gat) );
AND2XL U_g2115P1229 (.A(G3165P927gat), .B(G3167P931_bgat), .Y(G2115P1229gat) );
OR2XL U_g5330P1231 (.A(G3282P928gat), .B(G5322P932gat), .Y(G5330P1231gat) );
INVXL U_g5206P929_b (.A(G5206P929gat), .Y(G5206P929_bgat) );
OR2XL U_g5215P1233 (.A(G5209P925gat), .B(G5206P929_bgat), .Y(G5215P1233gat) );
OR2XL U_g3484P1241 (.A(G5178P934gat), .B(G2802P950_bgat), .Y(G3484P1241gat) );
AND3XL U_g3955P1242 (.A(G3897P935gat), .B(G3906P938gat), .C(G3915P941gat), .Y(G3955P1242gat) );
INVXL U_g3897P935_b (.A(G3897P935gat), .Y(G3897P935_bgat) );
INVXL U_g3906P938_b (.A(G3906P938gat), .Y(G3906P938_bgat) );
AND3XL U_g3958P1243 (.A(G3897P935_bgat), .B(G3906P938_bgat), .C(G3915P941gat), .Y(G3958P1243gat) );
INVXL U_g5396P1110_b (.A(G5396P1110gat), .Y(G5396P1110_bgat) );
OR2XL U_g5405P1264 (.A(G5399P946gat), .B(G5396P1110_bgat), .Y(G5405P1264gat) );
AND2XL U_g1875P1279 (.A(G54P20gat), .B(G3137P914_bgat), .Y(G1875P1279gat) );
AND3XL U_g4067P1284 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3012P1132gat), .Y(G4067P1284gat) );
AND3XL U_g4070P1285 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2942P1137gat), .Y(G4070P1285gat) );
AND3XL U_g4073P1286 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2939P1144gat), .Y(G4073P1286gat) );
AND3XL U_g4009P1287 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2623P1167gat), .Y(G4009P1287gat) );
AND3XL U_g4012P1288 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2619P1171gat), .Y(G4012P1288gat) );
AND3XL U_g4015P1289 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2615P1155gat), .Y(G4015P1289gat) );
AND3XL U_g4018P1290 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2611P1159gat), .Y(G4018P1290gat) );
AND3XL U_g3839P1291 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3021P1123gat), .Y(G3839P1291gat) );
AND3XL U_g3842P1292 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3018P1126gat), .Y(G3842P1292gat) );
AND3XL U_g3778P1293 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2717P1191gat), .Y(G3778P1293gat) );
AND3XL U_g3781P1294 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2713P1178gat), .Y(G3781P1294gat) );
AND3XL U_g3784P1295 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2709P1183gat), .Y(G3784P1295gat) );
AND3XL U_g3787P1296 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G2705P1186gat), .Y(G3787P1296gat) );
INVXL U_g534P149_b (.A(G534P149gat), .Y(G534P149_bgat) );
OR2XL U_g2066P1299 (.A(G534P149_bgat), .B(G3139P917gat), .Y(G2066P1299gat) );
OR2XL U_g1810P1300 (.A(G534P149_bgat), .B(G3139P917gat), .Y(G1810P1300gat) );
INVXL U_g523P148_b (.A(G523P148gat), .Y(G523P148_bgat) );
OR2XL U_g1792P1303 (.A(G523P148_bgat), .B(G3143P919gat), .Y(G1792P1303gat) );
OR2XL U_g2041P1304 (.A(G523P148_bgat), .B(G3143P919gat), .Y(G2041P1304gat) );
INVXL U_g5304P1133_b (.A(G5304P1133gat), .Y(G5304P1133_bgat) );
OR2XL U_g3891P1305 (.A(G5307P862gat), .B(G5304P1133_bgat), .Y(G3891P1305gat) );
INVXL U_g2019P978_b (.A(G2019P978gat), .Y(G2019P978_bgat) );
INVXL U_g2020P1130_b (.A(G2020P1130gat), .Y(G2020P1130_bgat) );
OR2XL U_g2021P1306 (.A(G2019P978_bgat), .B(G2020P1130_bgat), .Y(G2021P1306gat) );
INVXL U_g1777P979_b (.A(G1777P979gat), .Y(G1777P979_bgat) );
INVXL U_g1776P1131_b (.A(G1776P1131gat), .Y(G1776P1131_bgat) );
OR2XL U_g1778P1307 (.A(G1777P979_bgat), .B(G1776P1131_bgat), .Y(G1778P1307gat) );
INVXL U_g503P146_b (.A(G503P146gat), .Y(G503P146_bgat) );
OR2XL U_g2008P1310 (.A(G503P146_bgat), .B(G3151P923gat), .Y(G2008P1310gat) );
OR2XL U_g1765P1311 (.A(G503P146_bgat), .B(G3151P923gat), .Y(G1765P1311gat) );
OR2XL U_g2098P1314 (.A(G490P145_bgat), .B(G3155P924gat), .Y(G2098P1314gat) );
OR2XL U_g1756P1316 (.A(G490P145_bgat), .B(G3155P924gat), .Y(G1756P1316gat) );
INVXL U_g479P144_b (.A(G479P144gat), .Y(G479P144_bgat) );
OR2XL U_g1728P1320 (.A(G479P144_bgat), .B(G3161P926gat), .Y(G1728P1320gat) );
OR2XL U_g1983P1321 (.A(G479P144_bgat), .B(G3161P926gat), .Y(G1983P1321gat) );
INVXL U_g468P143_b (.A(G468P143gat), .Y(G468P143_bgat) );
OR2XL U_g1050P1324 (.A(G468P143_bgat), .B(G2794P947gat), .Y(G1050P1324gat) );
OR2XL U_g1306P1325 (.A(G468P143_bgat), .B(G2794P947gat), .Y(G1306P1325gat) );
INVXL U_g457P142_b (.A(G457P142gat), .Y(G457P142_bgat) );
OR2XL U_g1288P1328 (.A(G457P142_bgat), .B(G2798P948gat), .Y(G1288P1328gat) );
OR2XL U_g1032P1329 (.A(G457P142_bgat), .B(G2798P948gat), .Y(G1032P1329gat) );
INVXL U_g3338P1003_b (.A(G3338P1003gat), .Y(G3338P1003_bgat) );
AND2XL U_g3353P1330 (.A(G3347P1002gat), .B(G3338P1003_bgat), .Y(G3353P1330gat) );
INVXL U_g3331P1005_b (.A(G3331P1005gat), .Y(G3331P1005_bgat) );
AND2XL U_g3350P1331 (.A(G3343P1004gat), .B(G3331P1005_bgat), .Y(G3350P1331gat) );
INVXL U_g446P141_b (.A(G446P141gat), .Y(G446P141_bgat) );
OR2XL U_g1021P1332 (.A(G446P141_bgat), .B(G2802P950gat), .Y(G1021P1332gat) );
OR2XL U_g1277P1333 (.A(G446P141_bgat), .B(G2802P950gat), .Y(G1277P1333gat) );
INVXL U_g435P140_b (.A(G435P140gat), .Y(G435P140_bgat) );
OR2XL U_g1331P1336 (.A(G435P140_bgat), .B(G2784P944gat), .Y(G1331P1336gat) );
OR2XL U_g1087P1337 (.A(G435P140_bgat), .B(G2784P944gat), .Y(G1087P1337gat) );
OR2XL U_g1078P1340 (.A(G422P139_bgat), .B(G2788P945gat), .Y(G1078P1340gat) );
OR2XL U_g1421P1342 (.A(G422P139_bgat), .B(G2788P945gat), .Y(G1421P1342gat) );
INVXL U_g411P138_b (.A(G411P138gat), .Y(G411P138_bgat) );
OR2XL U_g1132P1346 (.A(G411P138_bgat), .B(G2772P937gat), .Y(G1132P1346gat) );
OR2XL U_g1389P1347 (.A(G411P138_bgat), .B(G2772P937gat), .Y(G1389P1347gat) );
INVXL U_g400P137_b (.A(G400P137gat), .Y(G400P137_bgat) );
OR2XL U_g1364P1350 (.A(G400P137_bgat), .B(G2776P939gat), .Y(G1364P1350gat) );
OR2XL U_g1114P1351 (.A(G400P137_bgat), .B(G2776P939gat), .Y(G1114P1351gat) );
INVXL U_g389P136_b (.A(G389P136gat), .Y(G389P136_bgat) );
OR2XL U_g1098P1354 (.A(G389P136_bgat), .B(G2780P940gat), .Y(G1098P1354gat) );
OR2XL U_g1343P1355 (.A(G389P136_bgat), .B(G2780P940gat), .Y(G1343P1355gat) );
OR2XL U_g1429P1358 (.A(G374P134_bgat), .B(G2767P936gat), .Y(G1429P1358gat) );
OR2XL U_g1150P1360 (.A(G374P134_bgat), .B(G2767P936gat), .Y(G1150P1360gat) );
INVXL U_g5126P912_b (.A(G5126P912gat), .Y(G5126P912_bgat) );
OR2XL U_g3453P1361 (.A(G5126P912_bgat), .B(G3137P914gat), .Y(G3453P1361gat) );
OR2XL U_g4756P1363 (.A(G3137P914gat), .B(G1875P1279gat), .Y(G4756P1363gat) );
OR2XL U_g3444P1368 (.A(G3139P917_bgat), .B(G3143P919gat), .Y(G3444P1368gat) );
OR2XL U_g3443P1369 (.A(G3139P917gat), .B(G3143P919_bgat), .Y(G3443P1369gat) );
OR2XL U_g3461P1370 (.A(G3147P723_bgat), .B(G3151P923gat), .Y(G3461P1370gat) );
INVXL U_g3517P1214_b (.A(G3517P1214gat), .Y(G3517P1214_bgat) );
INVXL U_g3516P1215_b (.A(G3516P1215gat), .Y(G3516P1215_bgat) );
AND2XL U_g3518P1371 (.A(G3517P1214_bgat), .B(G3516P1215_bgat), .Y(G3518P1371gat) );
INVXL U_g3514P1057_b (.A(G3514P1057gat), .Y(G3514P1057_bgat) );
INVXL U_g3513P1216_b (.A(G3513P1216gat), .Y(G3513P1216_bgat) );
AND2XL U_g3515P1372 (.A(G3514P1057_bgat), .B(G3513P1216_bgat), .Y(G3515P1372gat) );
OR2XL U_g5150P1373 (.A(G3155P924_bgat), .B(G3161P926gat), .Y(G5150P1373gat) );
INVXL U_g5214P1220_b (.A(G5214P1220gat), .Y(G5214P1220_bgat) );
INVXL U_g5215P1233_b (.A(G5215P1233gat), .Y(G5215P1233_bgat) );
OR2XL U_g5239P1374 (.A(G5214P1220_bgat), .B(G5215P1233_bgat), .Y(G5239P1374gat) );
OR2XL U_g5151P1375 (.A(G3155P924gat), .B(G3161P926_bgat), .Y(G5151P1375gat) );
OR2XL U_g5160P1380 (.A(G3165P927_bgat), .B(G3167P931gat), .Y(G5160P1380gat) );
OR2XL U_g5161P1385 (.A(G3165P927gat), .B(G3167P931_bgat), .Y(G5161P1385gat) );
INVXL U_g3282P928_b (.A(G3282P928gat), .Y(G3282P928_bgat) );
INVXL U_g5322P932_b (.A(G5322P932gat), .Y(G5322P932_bgat) );
OR2XL U_g5331P1387 (.A(G3282P928_bgat), .B(G5322P932_bgat), .Y(G5331P1387gat) );
INVXL U_g5178P934_b (.A(G5178P934gat), .Y(G5178P934_bgat) );
OR2XL U_g3485P1388 (.A(G5178P934_bgat), .B(G2802P950gat), .Y(G3485P1388gat) );
INVXL U_g3915P941_b (.A(G3915P941gat), .Y(G3915P941_bgat) );
AND3XL U_g3957P1389 (.A(G3897P935gat), .B(G3906P938_bgat), .C(G3915P941_bgat), .Y(G3957P1389gat) );
OR2XL U_g5194P1390 (.A(G2767P936_bgat), .B(G2772P937gat), .Y(G5194P1390gat) );
OR2XL U_g5195P1391 (.A(G2767P936gat), .B(G2772P937_bgat), .Y(G5195P1391gat) );
AND3XL U_g3954P1392 (.A(G3897P935_bgat), .B(G3906P938gat), .C(G3915P941_bgat), .Y(G3954P1392gat) );
OR2XL U_g5204P1393 (.A(G2776P939_bgat), .B(G2780P940gat), .Y(G5204P1393gat) );
OR2XL U_g5205P1394 (.A(G2776P939gat), .B(G2780P940_bgat), .Y(G5205P1394gat) );
OR2XL U_g3466P1395 (.A(G2784P944_bgat), .B(G2788P945gat), .Y(G3466P1395gat) );
OR2XL U_g3467P1396 (.A(G2784P944gat), .B(G2788P945_bgat), .Y(G3467P1396gat) );
INVXL U_g5399P946_b (.A(G5399P946gat), .Y(G5399P946_bgat) );
OR2XL U_g5404P1397 (.A(G5399P946_bgat), .B(G5396P1110gat), .Y(G5404P1397gat) );
OR2XL U_g3475P1398 (.A(G2794P947_bgat), .B(G2798P948gat), .Y(G3475P1398gat) );
OR2XL U_g3476P1399 (.A(G2794P947gat), .B(G2798P948_bgat), .Y(G3476P1399gat) );
OR2XL U_g1876P1400 (.A(G54P20gat), .B(G3137P914gat), .Y(G1876P1400gat) );
AND3XL U_g4021P1401 (.A(G4091P175_bgat), .B(G4092P176_bgat), .C(G3353P1330gat), .Y(G4021P1401gat) );
INVXL U_g5299P1122_b (.A(G5299P1122gat), .Y(G5299P1122_bgat) );
OR2XL U_g3881P1402 (.A(G5299P1122_bgat), .B(G5296P1127gat), .Y(G3881P1402gat) );
INVXL U_g2065P1124_b (.A(G2065P1124gat), .Y(G2065P1124_bgat) );
INVXL U_g2066P1299_b (.A(G2066P1299gat), .Y(G2066P1299_bgat) );
OR2XL U_g2067P1403 (.A(G2065P1124_bgat), .B(G2066P1299_bgat), .Y(G2067P1403gat) );
INVXL U_g1811P1125_b (.A(G1811P1125gat), .Y(G1811P1125_bgat) );
INVXL U_g1810P1300_b (.A(G1810P1300gat), .Y(G1810P1300_bgat) );
OR2XL U_g1812P1404 (.A(G1811P1125_bgat), .B(G1810P1300_bgat), .Y(G1812P1404gat) );
INVXL U_g5296P1127_b (.A(G5296P1127gat), .Y(G5296P1127_bgat) );
OR2XL U_g3882P1405 (.A(G5299P1122gat), .B(G5296P1127_bgat), .Y(G3882P1405gat) );
INVXL U_g1793P1128_b (.A(G1793P1128gat), .Y(G1793P1128_bgat) );
INVXL U_g1792P1303_b (.A(G1792P1303gat), .Y(G1792P1303_bgat) );
OR2XL U_g1794P1406 (.A(G1793P1128_bgat), .B(G1792P1303_bgat), .Y(G1794P1406gat) );
AND2XL U_g1866P1407 (.A(G1806P974gat), .B(G1778P1307gat), .Y(G1866P1407gat) );
INVXL U_g2040P1129_b (.A(G2040P1129gat), .Y(G2040P1129_bgat) );
INVXL U_g2041P1304_b (.A(G2041P1304gat), .Y(G2041P1304_bgat) );
OR2XL U_g2042P1408 (.A(G2040P1129_bgat), .B(G2041P1304_bgat), .Y(G2042P1408gat) );
AND2XL U_g2146P1409 (.A(G2059P975gat), .B(G2021P1306gat), .Y(G2146P1409gat) );
AND2XL U_g2142P1410 (.A(G2059P975gat), .B(G2021P1306gat), .Y(G2142P1410gat) );
INVXL U_g5307P862_b (.A(G5307P862gat), .Y(G5307P862_bgat) );
OR2XL U_g3890P1411 (.A(G5307P862_bgat), .B(G5304P1133gat), .Y(G3890P1411gat) );
INVXL U_g2007P1134_b (.A(G2007P1134gat), .Y(G2007P1134_bgat) );
INVXL U_g2008P1310_b (.A(G2008P1310gat), .Y(G2008P1310_bgat) );
OR2XL U_g2009P1416 (.A(G2007P1134_bgat), .B(G2008P1310_bgat), .Y(G2009P1416gat) );
INVXL U_g1766P1135_b (.A(G1766P1135gat), .Y(G1766P1135_bgat) );
INVXL U_g1765P1311_b (.A(G1765P1311gat), .Y(G1765P1311_bgat) );
OR2XL U_g1767P1417 (.A(G1766P1135_bgat), .B(G1765P1311_bgat), .Y(G1767P1417gat) );
INVXL U_g5315P1136_b (.A(G5315P1136gat), .Y(G5315P1136_bgat) );
OR2XL U_g5320P1418 (.A(G5315P1136_bgat), .B(G5312P1145gat), .Y(G5320P1418gat) );
INVXL U_g2097P1138_b (.A(G2097P1138gat), .Y(G2097P1138_bgat) );
INVXL U_g2098P1314_b (.A(G2098P1314gat), .Y(G2098P1314_bgat) );
OR2XL U_g2099P1419 (.A(G2097P1138_bgat), .B(G2098P1314_bgat), .Y(G2099P1419gat) );
INVXL U_g1757P1141_b (.A(G1757P1141gat), .Y(G1757P1141_bgat) );
INVXL U_g1756P1316_b (.A(G1756P1316gat), .Y(G1756P1316_bgat) );
OR2XL U_g1758P1420 (.A(G1757P1141_bgat), .B(G1756P1316_bgat), .Y(G1758P1420gat) );
INVXL U_g5312P1145_b (.A(G5312P1145gat), .Y(G5312P1145_bgat) );
OR2XL U_g5321P1421 (.A(G5315P1136gat), .B(G5312P1145_bgat), .Y(G5321P1421gat) );
INVXL U_g1729P1146_b (.A(G1729P1146gat), .Y(G1729P1146_bgat) );
INVXL U_g1728P1320_b (.A(G1728P1320gat), .Y(G1728P1320_bgat) );
OR2XL U_g1730P1422 (.A(G1729P1146_bgat), .B(G1728P1320_bgat), .Y(G1730P1422gat) );
INVXL U_g1982P1150_b (.A(G1982P1150gat), .Y(G1982P1150_bgat) );
INVXL U_g1983P1321_b (.A(G1983P1321gat), .Y(G1983P1321_bgat) );
OR2XL U_g1984P1423 (.A(G1982P1150_bgat), .B(G1983P1321_bgat), .Y(G1984P1423gat) );
INVXL U_g5276P1154_b (.A(G5276P1154gat), .Y(G5276P1154_bgat) );
OR2XL U_g5285P1424 (.A(G5276P1154_bgat), .B(G5279P1170gat), .Y(G5285P1424gat) );
INVXL U_g1051P1156_b (.A(G1051P1156gat), .Y(G1051P1156_bgat) );
INVXL U_g1050P1324_b (.A(G1050P1324gat), .Y(G1050P1324_bgat) );
OR2XL U_g1052P1426 (.A(G1051P1156_bgat), .B(G1050P1324_bgat), .Y(G1052P1426gat) );
INVXL U_g1305P1157_b (.A(G1305P1157gat), .Y(G1305P1157_bgat) );
INVXL U_g1306P1325_b (.A(G1306P1325gat), .Y(G1306P1325_bgat) );
OR2XL U_g1307P1427 (.A(G1305P1157_bgat), .B(G1306P1325_bgat), .Y(G1307P1427gat) );
INVXL U_g1287P1160_b (.A(G1287P1160gat), .Y(G1287P1160_bgat) );
INVXL U_g1288P1328_b (.A(G1288P1328gat), .Y(G1288P1328_bgat) );
OR2XL U_g1289P1428 (.A(G1287P1160_bgat), .B(G1288P1328_bgat), .Y(G1289P1428gat) );
INVXL U_g1033P1161_b (.A(G1033P1161gat), .Y(G1033P1161_bgat) );
INVXL U_g1032P1329_b (.A(G1032P1329gat), .Y(G1032P1329_bgat) );
OR2XL U_g1034P1429 (.A(G1033P1161_bgat), .B(G1032P1329_bgat), .Y(G1034P1429gat) );
INVXL U_g1022P1164_b (.A(G1022P1164gat), .Y(G1022P1164_bgat) );
INVXL U_g1021P1332_b (.A(G1021P1332gat), .Y(G1021P1332_bgat) );
OR2XL U_g1023P1432 (.A(G1022P1164_bgat), .B(G1021P1332_bgat), .Y(G1023P1432gat) );
INVXL U_g1276P1165_b (.A(G1276P1165gat), .Y(G1276P1165_bgat) );
INVXL U_g1277P1333_b (.A(G1277P1333gat), .Y(G1277P1333_bgat) );
OR2XL U_g1278P1433 (.A(G1276P1165_bgat), .B(G1277P1333_bgat), .Y(G1278P1433gat) );
INVXL U_g5268P1166_b (.A(G5268P1166gat), .Y(G5268P1166_bgat) );
OR2XL U_g3870P1434 (.A(G5268P1166_bgat), .B(G5271P1187gat), .Y(G3870P1434gat) );
INVXL U_g1330P1168_b (.A(G1330P1168gat), .Y(G1330P1168_bgat) );
INVXL U_g1331P1336_b (.A(G1331P1336gat), .Y(G1331P1336_bgat) );
OR2XL U_g1332P1435 (.A(G1330P1168_bgat), .B(G1331P1336_bgat), .Y(G1332P1435gat) );
INVXL U_g1088P1169_b (.A(G1088P1169gat), .Y(G1088P1169_bgat) );
INVXL U_g1087P1337_b (.A(G1087P1337gat), .Y(G1087P1337_bgat) );
OR2XL U_g1089P1436 (.A(G1088P1169_bgat), .B(G1087P1337_bgat), .Y(G1089P1436gat) );
INVXL U_g5279P1170_b (.A(G5279P1170gat), .Y(G5279P1170_bgat) );
OR2XL U_g5284P1437 (.A(G5276P1154gat), .B(G5279P1170_bgat), .Y(G5284P1437gat) );
INVXL U_g1079P1172_b (.A(G1079P1172gat), .Y(G1079P1172_bgat) );
INVXL U_g1078P1340_b (.A(G1078P1340gat), .Y(G1078P1340_bgat) );
OR2XL U_g1080P1438 (.A(G1079P1172_bgat), .B(G1078P1340_bgat), .Y(G1080P1438gat) );
INVXL U_g1420P1175_b (.A(G1420P1175gat), .Y(G1420P1175_bgat) );
INVXL U_g1421P1342_b (.A(G1421P1342gat), .Y(G1421P1342_bgat) );
OR2XL U_g1422P1439 (.A(G1420P1175_bgat), .B(G1421P1342_bgat), .Y(G1422P1439gat) );
INVXL U_g5263P1179_b (.A(G5263P1179gat), .Y(G5263P1179_bgat) );
OR2XL U_g3860P1441 (.A(G5263P1179_bgat), .B(G5260P1182gat), .Y(G3860P1441gat) );
INVXL U_g1133P1180_b (.A(G1133P1180gat), .Y(G1133P1180_bgat) );
INVXL U_g1132P1346_b (.A(G1132P1346gat), .Y(G1132P1346_bgat) );
OR2XL U_g1134P1442 (.A(G1133P1180_bgat), .B(G1132P1346_bgat), .Y(G1134P1442gat) );
INVXL U_g1388P1181_b (.A(G1388P1181gat), .Y(G1388P1181_bgat) );
INVXL U_g1389P1347_b (.A(G1389P1347gat), .Y(G1389P1347_bgat) );
OR2XL U_g1390P1443 (.A(G1388P1181_bgat), .B(G1389P1347_bgat), .Y(G1390P1443gat) );
INVXL U_g5260P1182_b (.A(G5260P1182gat), .Y(G5260P1182_bgat) );
OR2XL U_g3861P1444 (.A(G5263P1179gat), .B(G5260P1182_bgat), .Y(G3861P1444gat) );
INVXL U_g1363P1184_b (.A(G1363P1184gat), .Y(G1363P1184_bgat) );
INVXL U_g1364P1350_b (.A(G1364P1350gat), .Y(G1364P1350_bgat) );
OR2XL U_g1365P1445 (.A(G1363P1184_bgat), .B(G1364P1350_bgat), .Y(G1365P1445gat) );
INVXL U_g1115P1185_b (.A(G1115P1185gat), .Y(G1115P1185_bgat) );
INVXL U_g1114P1351_b (.A(G1114P1351gat), .Y(G1114P1351_bgat) );
OR2XL U_g1116P1446 (.A(G1115P1185_bgat), .B(G1114P1351_bgat), .Y(G1116P1446gat) );
INVXL U_g5271P1187_b (.A(G5271P1187gat), .Y(G5271P1187_bgat) );
OR2XL U_g3869P1447 (.A(G5268P1166gat), .B(G5271P1187_bgat), .Y(G3869P1447gat) );
INVXL U_g1099P1188_b (.A(G1099P1188gat), .Y(G1099P1188_bgat) );
INVXL U_g1098P1354_b (.A(G1098P1354gat), .Y(G1098P1354_bgat) );
OR2XL U_g1100P1448 (.A(G1099P1188_bgat), .B(G1098P1354_bgat), .Y(G1100P1448gat) );
INVXL U_g1342P1189_b (.A(G1342P1189gat), .Y(G1342P1189_bgat) );
INVXL U_g1343P1355_b (.A(G1343P1355gat), .Y(G1343P1355_bgat) );
OR2XL U_g1344P1449 (.A(G1342P1189_bgat), .B(G1343P1355_bgat), .Y(G1344P1449gat) );
INVXL U_g1428P1192_b (.A(G1428P1192gat), .Y(G1428P1192_bgat) );
INVXL U_g1429P1358_b (.A(G1429P1358gat), .Y(G1429P1358_bgat) );
OR2XL U_g1430P1451 (.A(G1428P1192_bgat), .B(G1429P1358_bgat), .Y(G1430P1451gat) );
INVXL U_g1151P1195_b (.A(G1151P1195gat), .Y(G1151P1195_bgat) );
INVXL U_g1150P1360_b (.A(G1150P1360gat), .Y(G1150P1360_bgat) );
OR2XL U_g1152P1452 (.A(G1151P1195_bgat), .B(G1150P1360_bgat), .Y(G1152P1452gat) );
INVXL U_g3452P1196_b (.A(G3452P1196gat), .Y(G3452P1196_bgat) );
INVXL U_g3453P1361_b (.A(G3453P1361gat), .Y(G3453P1361_bgat) );
OR2XL U_g3454P1453 (.A(G3452P1196_bgat), .B(G3453P1361_bgat), .Y(G3454P1453gat) );
INVXL U_g3444P1368_b (.A(G3444P1368gat), .Y(G3444P1368_bgat) );
INVXL U_g3443P1369_b (.A(G3443P1369gat), .Y(G3443P1369_bgat) );
OR2XL U_g3445P1455 (.A(G3444P1368_bgat), .B(G3443P1369_bgat), .Y(G3445P1455gat) );
INVXL U_g3462P1210_b (.A(G3462P1210gat), .Y(G3462P1210_bgat) );
INVXL U_g3461P1370_b (.A(G3461P1370gat), .Y(G3461P1370_bgat) );
OR2XL U_g3463P1456 (.A(G3462P1210_bgat), .B(G3461P1370_bgat), .Y(G3463P1456gat) );
INVXL U_g3518P1371_b (.A(G3518P1371gat), .Y(G3518P1371_bgat) );
INVXL U_g3515P1372_b (.A(G3515P1372gat), .Y(G3515P1372_bgat) );
OR2XL U_g5236P1457 (.A(G3518P1371_bgat), .B(G3515P1372_bgat), .Y(G5236P1457gat) );
INVXL U_g5150P1373_b (.A(G5150P1373gat), .Y(G5150P1373_bgat) );
INVXL U_g5151P1375_b (.A(G5151P1375gat), .Y(G5151P1375_bgat) );
OR2XL U_g5219P1458 (.A(G5150P1373_bgat), .B(G5151P1375_bgat), .Y(G5219P1458gat) );
INVXL U_g5160P1380_b (.A(G5160P1380gat), .Y(G5160P1380_bgat) );
INVXL U_g5161P1385_b (.A(G5161P1385gat), .Y(G5161P1385_bgat) );
OR2XL U_g5216P1460 (.A(G5160P1380_bgat), .B(G5161P1385_bgat), .Y(G5216P1460gat) );
INVXL U_g5330P1231_b (.A(G5330P1231gat), .Y(G5330P1231_bgat) );
INVXL U_g5331P1387_b (.A(G5331P1387gat), .Y(G5331P1387_bgat) );
OR2XL U_g5386P1461 (.A(G5330P1231_bgat), .B(G5331P1387_bgat), .Y(G5386P1461gat) );
INVXL U_g3484P1241_b (.A(G3484P1241gat), .Y(G3484P1241_bgat) );
INVXL U_g3485P1388_b (.A(G3485P1388gat), .Y(G3485P1388_bgat) );
OR2XL U_g3486P1464 (.A(G3484P1241_bgat), .B(G3485P1388_bgat), .Y(G3486P1464gat) );
INVXL U_g3955P1242_b (.A(G3955P1242gat), .Y(G3955P1242_bgat) );
INVXL U_g3954P1392_b (.A(G3954P1392gat), .Y(G3954P1392_bgat) );
AND2XL U_g3956P1465 (.A(G3955P1242_bgat), .B(G3954P1392_bgat), .Y(G3956P1465gat) );
INVXL U_g3958P1243_b (.A(G3958P1243gat), .Y(G3958P1243_bgat) );
INVXL U_g3957P1389_b (.A(G3957P1389gat), .Y(G3957P1389_bgat) );
AND2XL U_g3959P1466 (.A(G3958P1243_bgat), .B(G3957P1389_bgat), .Y(G3959P1466gat) );
INVXL U_g5194P1390_b (.A(G5194P1390gat), .Y(G5194P1390_bgat) );
INVXL U_g5195P1391_b (.A(G5195P1391gat), .Y(G5195P1391_bgat) );
OR2XL U_g5229P1467 (.A(G5194P1390_bgat), .B(G5195P1391_bgat), .Y(G5229P1467gat) );
INVXL U_g5204P1393_b (.A(G5204P1393gat), .Y(G5204P1393_bgat) );
INVXL U_g5205P1394_b (.A(G5205P1394gat), .Y(G5205P1394_bgat) );
OR2XL U_g5226P1468 (.A(G5204P1393_bgat), .B(G5205P1394_bgat), .Y(G5226P1468gat) );
INVXL U_g3466P1395_b (.A(G3466P1395gat), .Y(G3466P1395_bgat) );
INVXL U_g3467P1396_b (.A(G3467P1396gat), .Y(G3467P1396_bgat) );
OR2XL U_g3468P1469 (.A(G3466P1395_bgat), .B(G3467P1396_bgat), .Y(G3468P1469gat) );
INVXL U_g5405P1264_b (.A(G5405P1264gat), .Y(G5405P1264_bgat) );
INVXL U_g5404P1397_b (.A(G5404P1397gat), .Y(G5404P1397_bgat) );
OR2XL U_g5425P1470 (.A(G5405P1264_bgat), .B(G5404P1397_bgat), .Y(G5425P1470gat) );
INVXL U_g3475P1398_b (.A(G3475P1398gat), .Y(G3475P1398_bgat) );
INVXL U_g3476P1399_b (.A(G3476P1399gat), .Y(G3476P1399_bgat) );
OR2XL U_g3477P1471 (.A(G3475P1398_bgat), .B(G3476P1399_bgat), .Y(G3477P1471gat) );
INVXL U_g54P20_b (.A(G54P20gat), .Y(G54P20_bgat) );
OR2XL U_g1877P1472 (.A(G54P20_bgat), .B(G3137P914_bgat), .Y(G1877P1472gat) );
INVXL U_g3881P1402_b (.A(G3881P1402gat), .Y(G3881P1402_bgat) );
INVXL U_g3882P1405_b (.A(G3882P1405gat), .Y(G3882P1405_bgat) );
OR2XL U_g3883P1473 (.A(G3881P1402_bgat), .B(G3882P1405_bgat), .Y(G3883P1473gat) );
AND3XL U_g2147P1476 (.A(G2081P970gat), .B(G2021P1306gat), .C(G2042P1408gat), .Y(G2147P1476gat) );
AND3XL U_g2143P1477 (.A(G2081P970gat), .B(G2021P1306gat), .C(G2042P1408gat), .Y(G2143P1477gat) );
AND4XL U_g2133P1478 (.A(G2081P970gat), .B(G2021P1306gat), .C(G2042P1408gat), .D(G2009P1416gat), .Y(G2133P1478gat) );
AND2XL U_g2152P1479 (.A(G2081P970gat), .B(G2042P1408gat), .Y(G2152P1479gat) );
AND2XL U_g2149P1480 (.A(G2081P970gat), .B(G2042P1408gat), .Y(G2149P1480gat) );
AND3XL U_g1867P1481 (.A(G1823P971gat), .B(G1778P1307gat), .C(G1794P1406gat), .Y(G1867P1481gat) );
AND4XL U_g1861P1482 (.A(G1823P971gat), .B(G1778P1307gat), .C(G1794P1406gat), .D(G1767P1417gat), .Y(G1861P1482gat) );
AND2XL U_g1870P1483 (.A(G1823P971gat), .B(G1794P1406gat), .Y(G1870P1483gat) );
AND3XL U_g1860P1486 (.A(G1806P974gat), .B(G1778P1307gat), .C(G1767P1417gat), .Y(G1860P1486gat) );
AND3XL U_g2132P1489 (.A(G2059P975gat), .B(G2021P1306gat), .C(G2009P1416gat), .Y(G2132P1489gat) );
INVXL U_g3891P1305_b (.A(G3891P1305gat), .Y(G3891P1305_bgat) );
INVXL U_g3890P1411_b (.A(G3890P1411gat), .Y(G3890P1411_bgat) );
OR2XL U_g3892P1490 (.A(G3891P1305_bgat), .B(G3890P1411_bgat), .Y(G3892P1490gat) );
AND2XL U_g2131P1493 (.A(G2036P864gat), .B(G2009P1416gat), .Y(G2131P1493gat) );
AND2XL U_g1859P1495 (.A(G1789P865gat), .B(G1767P1417gat), .Y(G1859P1495gat) );
INVXL U_g5320P1418_b (.A(G5320P1418gat), .Y(G5320P1418_bgat) );
INVXL U_g5321P1421_b (.A(G5321P1421gat), .Y(G5321P1421_bgat) );
OR2XL U_g5389P1499 (.A(G5320P1418_bgat), .B(G5321P1421_bgat), .Y(G5389P1499gat) );
AND2XL U_g2158P1501 (.A(G2099P1419gat), .B(G1984P1423gat), .Y(G2158P1501gat) );
AND3XL U_g2120P1503 (.A(G3165P927_bgat), .B(G2001P987gat), .C(G1984P1423gat), .Y(G2120P1503gat) );
AND4XL U_g2117P1504 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G2001P987gat), .D(G1984P1423gat), .Y(G2117P1504gat) );
AND3XL U_g2123P1505 (.A(G3165P927_bgat), .B(G2001P987gat), .C(G1984P1423gat), .Y(G2123P1505gat) );
AND2XL U_g2124P1506 (.A(G2001P987gat), .B(G1984P1423gat), .Y(G2124P1506gat) );
AND2XL U_g1855P1507 (.A(G1758P1420gat), .B(G1730P1422gat), .Y(G1855P1507gat) );
AND4XL U_g1847P1509 (.A(G3165P927_bgat), .B(G3167P931_bgat), .C(G1749P988gat), .D(G1730P1422gat), .Y(G1847P1509gat) );
AND3XL U_g1853P1510 (.A(G3165P927_bgat), .B(G1749P988gat), .C(G1730P1422gat), .Y(G1853P1510gat) );
AND3XL U_g1850P1511 (.A(G3165P927_bgat), .B(G1749P988gat), .C(G1730P1422gat), .Y(G1850P1511gat) );
AND2XL U_g1854P1512 (.A(G1749P988gat), .B(G1730P1422gat), .Y(G1854P1512gat) );
AND2XL U_g1856P1513 (.A(G1749P988gat), .B(G1730P1422gat), .Y(G1856P1513gat) );
INVXL U_g5285P1424_b (.A(G5285P1424gat), .Y(G5285P1424_bgat) );
INVXL U_g5284P1437_b (.A(G5284P1437gat), .Y(G5284P1437_bgat) );
OR2XL U_g5379P1518 (.A(G5285P1424_bgat), .B(G5284P1437_bgat), .Y(G5379P1518gat) );
AND3XL U_g1173P1523 (.A(G1052P1426gat), .B(G1034P1429gat), .C(G1080P1438gat), .Y(G1173P1523gat) );
AND2XL U_g1177P1524 (.A(G1052P1426gat), .B(G1080P1438gat), .Y(G1177P1524gat) );
AND3XL U_g1169P1525 (.A(G1064P996gat), .B(G1034P1429gat), .C(G1023P1432gat), .Y(G1169P1525gat) );
AND2XL U_g1171P1526 (.A(G1064P996gat), .B(G1034P1429gat), .Y(G1171P1526gat) );
AND2XL U_g1174P1527 (.A(G1064P996gat), .B(G1034P1429gat), .Y(G1174P1527gat) );
AND2XL U_g1481P1528 (.A(G1307P1427gat), .B(G1422P1439gat), .Y(G1481P1528gat) );
AND3XL U_g1444P1531 (.A(G1307P1427gat), .B(G1289P1428gat), .C(G1422P1439gat), .Y(G1444P1531gat) );
AND2XL U_g1445P1533 (.A(G1318P997gat), .B(G1289P1428gat), .Y(G1445P1533gat) );
AND3XL U_g1440P1534 (.A(G1318P997gat), .B(G1289P1428gat), .C(G1278P1433gat), .Y(G1440P1534gat) );
AND2XL U_g1442P1535 (.A(G1318P997gat), .B(G1289P1428gat), .Y(G1442P1535gat) );
OR2XL U_g5295P1536 (.A(G5289P1158gat), .B(G3350P1331_bgat), .Y(G5295P1536gat) );
AND2XL U_g1439P1539 (.A(G1301P1000gat), .B(G1278P1433gat), .Y(G1439P1539gat) );
AND2XL U_g1168P1542 (.A(G1046P1001gat), .B(G1023P1432gat), .Y(G1168P1542gat) );
INVXL U_g3870P1434_b (.A(G3870P1434gat), .Y(G3870P1434_bgat) );
INVXL U_g3869P1447_b (.A(G3869P1447gat), .Y(G3869P1447_bgat) );
OR2XL U_g3871P1548 (.A(G3870P1434_bgat), .B(G3869P1447_bgat), .Y(G3871P1548gat) );
AND4XL U_g1170P1555 (.A(G1071P1014gat), .B(G1052P1426gat), .C(G1034P1429gat), .D(G1023P1432gat), .Y(G1170P1555gat) );
AND3XL U_g1175P1556 (.A(G1071P1014gat), .B(G1052P1426gat), .C(G1034P1429gat), .Y(G1175P1556gat) );
AND3XL U_g1172P1557 (.A(G1071P1014gat), .B(G1052P1426gat), .C(G1034P1429gat), .Y(G1172P1557gat) );
AND2XL U_g1176P1558 (.A(G1071P1014gat), .B(G1052P1426gat), .Y(G1176P1558gat) );
AND2XL U_g1178P1559 (.A(G1071P1014gat), .B(G1052P1426gat), .Y(G1178P1559gat) );
AND3XL U_g1443P1562 (.A(G1324P1017gat), .B(G1307P1427gat), .C(G1289P1428gat), .Y(G1443P1562gat) );
AND4XL U_g1441P1563 (.A(G1324P1017gat), .B(G1307P1427gat), .C(G1289P1428gat), .D(G1278P1433gat), .Y(G1441P1563gat) );
AND3XL U_g1446P1564 (.A(G1324P1017gat), .B(G1307P1427gat), .C(G1289P1428gat), .Y(G1446P1564gat) );
AND2XL U_g1447P1565 (.A(G1324P1017gat), .B(G1307P1427gat), .Y(G1447P1565gat) );
INVXL U_g3860P1441_b (.A(G3860P1441gat), .Y(G3860P1441_bgat) );
INVXL U_g3861P1444_b (.A(G3861P1444gat), .Y(G3861P1444_bgat) );
OR2XL U_g3862P1566 (.A(G3860P1441_bgat), .B(G3861P1444_bgat), .Y(G3862P1566gat) );
AND3XL U_g1189P1567 (.A(G1145P1020gat), .B(G1116P1446gat), .C(G1100P1448gat), .Y(G1189P1567gat) );
AND4XL U_g1183P1568 (.A(G1145P1020gat), .B(G1089P1436gat), .C(G1116P1446gat), .D(G1100P1448gat), .Y(G1183P1568gat) );
AND2XL U_g1192P1569 (.A(G1145P1020gat), .B(G1116P1446gat), .Y(G1192P1569gat) );
AND4XL U_g1468P1572 (.A(G1390P1443gat), .B(G1365P1445gat), .C(G1344P1449gat), .D(G1430P1451gat), .Y(G1468P1572gat) );
AND3XL U_g1474P1573 (.A(G1390P1443gat), .B(G1365P1445gat), .C(G1430P1451gat), .Y(G1474P1573gat) );
AND2XL U_g1482P1575 (.A(G1390P1443gat), .B(G1430P1451gat), .Y(G1482P1575gat) );
AND3XL U_g1470P1576 (.A(G1404P1021gat), .B(G1365P1445gat), .C(G1344P1449gat), .Y(G1470P1576gat) );
AND3XL U_g1466P1577 (.A(G1404P1021gat), .B(G1365P1445gat), .C(G1344P1449gat), .Y(G1466P1577gat) );
AND4XL U_g1456P1578 (.A(G1404P1021gat), .B(G1332P1435gat), .C(G1365P1445gat), .D(G1344P1449gat), .Y(G1456P1578gat) );
AND2XL U_g1475P1579 (.A(G1404P1021gat), .B(G1365P1445gat), .Y(G1475P1579gat) );
AND2XL U_g1472P1580 (.A(G1404P1021gat), .B(G1365P1445gat), .Y(G1472P1580gat) );
AND2XL U_g1469P1583 (.A(G1382P1024gat), .B(G1344P1449gat), .Y(G1469P1583gat) );
AND2XL U_g1465P1584 (.A(G1382P1024gat), .B(G1344P1449gat), .Y(G1465P1584gat) );
AND3XL U_g1455P1585 (.A(G1382P1024gat), .B(G1332P1435gat), .C(G1344P1449gat), .Y(G1455P1585gat) );
AND2XL U_g1188P1587 (.A(G1128P1025gat), .B(G1100P1448gat), .Y(G1188P1587gat) );
AND3XL U_g1182P1588 (.A(G1128P1025gat), .B(G1089P1436gat), .C(G1100P1448gat), .Y(G1182P1588gat) );
AND2XL U_g1181P1590 (.A(G1111P1028gat), .B(G1089P1436gat), .Y(G1181P1590gat) );
AND2XL U_g1454P1593 (.A(G1359P1029gat), .B(G1332P1435gat), .Y(G1454P1593gat) );
AND4XL U_g1467P1596 (.A(G1412P1033gat), .B(G1390P1443gat), .C(G1365P1445gat), .D(G1344P1449gat), .Y(G1467P1596gat) );
AND5XL U_g1457P1597 (.A(G1412P1033gat), .B(G1332P1435gat), .C(G1390P1443gat), .D(G1365P1445gat), .E(G1344P1449gat), .Y(G1457P1597gat) );
AND4XL U_g1471P1598 (.A(G1412P1033gat), .B(G1390P1443gat), .C(G1365P1445gat), .D(G1344P1449gat), .Y(G1471P1598gat) );
AND3XL U_g1473P1599 (.A(G1412P1033gat), .B(G1390P1443gat), .C(G1365P1445gat), .Y(G1473P1599gat) );
AND2XL U_g1477P1600 (.A(G1412P1033gat), .B(G1390P1443gat), .Y(G1477P1600gat) );
AND3XL U_g1476P1601 (.A(G1412P1033gat), .B(G1390P1443gat), .C(G1365P1445gat), .Y(G1476P1601gat) );
AND4XL U_g1190P1603 (.A(G1160P1034gat), .B(G1134P1442gat), .C(G1116P1446gat), .D(G1100P1448gat), .Y(G1190P1603gat) );
AND5XL U_g1184P1604 (.A(G1160P1034gat), .B(G1089P1436gat), .C(G1134P1442gat), .D(G1116P1446gat), .E(G1100P1448gat), .Y(G1184P1604gat) );
AND2XL U_g1195P1605 (.A(G1160P1034gat), .B(G1134P1442gat), .Y(G1195P1605gat) );
AND3XL U_g1193P1606 (.A(G1160P1034gat), .B(G1134P1442gat), .C(G1116P1446gat), .Y(G1193P1606gat) );
AND4XL U_g1868P1609 (.A(G3137P914gat), .B(G1778P1307gat), .C(G1812P1404gat), .D(G1794P1406gat), .Y(G1868P1609gat) );
AND5XL U_g1862P1610 (.A(G3137P914gat), .B(G1778P1307gat), .C(G1812P1404gat), .D(G1794P1406gat), .E(G1767P1417gat), .Y(G1862P1610gat) );
AND2XL U_g1873P1611 (.A(G3137P914gat), .B(G1812P1404gat), .Y(G1873P1611gat) );
AND3XL U_g1871P1612 (.A(G3137P914gat), .B(G1812P1404gat), .C(G1794P1406gat), .Y(G1871P1612gat) );
AND4XL U_g2144P1613 (.A(G3137P914gat), .B(G2021P1306gat), .C(G2067P1403gat), .D(G2042P1408gat), .Y(G2144P1613gat) );
AND5XL U_g2134P1614 (.A(G3137P914gat), .B(G2021P1306gat), .C(G2067P1403gat), .D(G2042P1408gat), .E(G2009P1416gat), .Y(G2134P1614gat) );
AND4XL U_g2148P1615 (.A(G3137P914gat), .B(G2021P1306gat), .C(G2067P1403gat), .D(G2042P1408gat), .Y(G2148P1615gat) );
AND3XL U_g2150P1616 (.A(G3137P914gat), .B(G2067P1403gat), .C(G2042P1408gat), .Y(G2150P1616gat) );
AND2XL U_g2154P1617 (.A(G3137P914gat), .B(G2067P1403gat), .Y(G2154P1617gat) );
AND3XL U_g2153P1618 (.A(G3137P914gat), .B(G2067P1403gat), .C(G2042P1408gat), .Y(G2153P1618gat) );
AND4XL U_g2145P1620 (.A(G3137P914_bgat), .B(G2021P1306gat), .C(G2067P1403gat), .D(G2042P1408gat), .Y(G2145P1620gat) );
AND2XL U_g2159P1621 (.A(G3137P914_bgat), .B(G2067P1403gat), .Y(G2159P1621gat) );
AND3XL U_g2151P1622 (.A(G3137P914_bgat), .B(G2067P1403gat), .C(G2042P1408gat), .Y(G2151P1622gat) );
INVXL U_g5236P1457_b (.A(G5236P1457gat), .Y(G5236P1457_bgat) );
OR2XL U_g3532P1627 (.A(G5239P1374gat), .B(G5236P1457_bgat), .Y(G3532P1627gat) );
AND3XL U_g1851P1631 (.A(G3165P927_bgat), .B(G1758P1420gat), .C(G1730P1422gat), .Y(G1851P1631gat) );
AND3XL U_g2121P1633 (.A(G3165P927_bgat), .B(G2099P1419gat), .C(G1984P1423gat), .Y(G2121P1633gat) );
INVXL U_g3956P1465_b (.A(G3956P1465gat), .Y(G3956P1465_bgat) );
INVXL U_g3959P1466_b (.A(G3959P1466gat), .Y(G3959P1466_bgat) );
OR2XL U_g5422P1638 (.A(G3956P1465_bgat), .B(G3959P1466_bgat), .Y(G5422P1638gat) );
INVXL U_g132P60_b (.A(G132P60gat), .Y(G132P60_bgat) );
OR2XL U_g4107P1644 (.A(G132P60_bgat), .B(G3167P931gat), .Y(G4107P1644gat) );
AND5XL U_g1869P1645 (.A(G54P20gat), .B(G3137P914_bgat), .C(G1778P1307gat), .D(G1812P1404gat), .E(G1794P1406gat), .Y(G1869P1645gat) );
AND3XL U_g1874P1646 (.A(G54P20gat), .B(G3137P914_bgat), .C(G1812P1404gat), .Y(G1874P1646gat) );
INVXL U_g1876P1400_b (.A(G1876P1400gat), .Y(G1876P1400_bgat) );
INVXL U_g1877P1472_b (.A(G1877P1472gat), .Y(G1877P1472_bgat) );
OR2XL U_g1878P1647 (.A(G1876P1400_bgat), .B(G1877P1472_bgat), .Y(G1878P1647gat) );
AND4XL U_g1872P1648 (.A(G54P20gat), .B(G3137P914_bgat), .C(G1812P1404gat), .D(G1794P1406gat), .Y(G1872P1648gat) );
AND5XL U_g1191P1649 (.A(G4P1gat), .B(G1134P1442gat), .C(G1116P1446gat), .D(G1100P1448gat), .E(G1152P1452gat), .Y(G1191P1649gat) );
AND2XL U_g1197P1650 (.A(G4P1gat), .B(G1152P1452gat), .Y(G1197P1650gat) );
AND3XL U_g1196P1651 (.A(G4P1gat), .B(G1134P1442gat), .C(G1152P1452gat), .Y(G1196P1651gat) );
AND4XL U_g1194P1652 (.A(G4P1gat), .B(G1134P1442gat), .C(G1116P1446gat), .D(G1152P1452gat), .Y(G1194P1652gat) );
AND3XL U_g3837P1653 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1878P1647gat), .Y(G3837P1653gat) );
OR2XL U_g2155P1657 (.A(G2081P970gat), .B(G2154P1617gat), .Y(G2155P1657gat) );
OR3XL U_g4748P1658 (.A(G1823P971gat), .B(G1873P1611gat), .C(G1874P1646gat), .Y(G4748P1658gat) );
OR4XL U_g4740P1661 (.A(G1806P974gat), .B(G1870P1483gat), .C(G1871P1612gat), .D(G1872P1648gat), .Y(G4740P1661gat) );
INVXL U_g2059P975_b (.A(G2059P975gat), .Y(G2059P975_bgat) );
INVXL U_g2152P1479_b (.A(G2152P1479gat), .Y(G2152P1479_bgat) );
INVXL U_g2153P1618_b (.A(G2153P1618gat), .Y(G2153P1618_bgat) );
AND3XL U_g5009P1664 (.A(G2059P975_bgat), .B(G2152P1479_bgat), .C(G2153P1618_bgat), .Y(G5009P1664gat) );
OR4XL U_g4928P1665 (.A(G2059P975gat), .B(G2149P1480gat), .C(G2150P1616gat), .D(G2151P1622gat), .Y(G4928P1665gat) );
INVXL U_g2036P864_b (.A(G2036P864gat), .Y(G2036P864_bgat) );
INVXL U_g2146P1409_b (.A(G2146P1409gat), .Y(G2146P1409_bgat) );
INVXL U_g2147P1476_b (.A(G2147P1476gat), .Y(G2147P1476_bgat) );
INVXL U_g2148P1615_b (.A(G2148P1615gat), .Y(G2148P1615_bgat) );
AND4XL U_g5029P1668 (.A(G2036P864_bgat), .B(G2146P1409_bgat), .C(G2147P1476_bgat), .D(G2148P1615_bgat), .Y(G5029P1668gat) );
OR5XL U_g4941P1669 (.A(G2036P864gat), .B(G2142P1410gat), .C(G2143P1477gat), .D(G2144P1613gat), .E(G2145P1620gat), .Y(G4941P1669gat) );
OR5XL U_g4732P1670 (.A(G1789P865gat), .B(G1866P1407gat), .C(G1867P1481gat), .D(G1868P1609gat), .E(G1869P1645gat), .Y(G4732P1670gat) );
OR5XL U_g2135P1673 (.A(G2018P982gat), .B(G2133P1478gat), .C(G2132P1489gat), .D(G2131P1493gat), .E(G2134P1614gat), .Y(G2135P1673gat) );
OR5XL U_g1863P1675 (.A(G1775P983gat), .B(G1861P1482gat), .C(G1860P1486gat), .D(G1859P1495gat), .E(G1862P1610gat), .Y(G1863P1675gat) );
INVXL U_g5389P1499_b (.A(G5389P1499gat), .Y(G5389P1499_bgat) );
OR2XL U_g5394P1676 (.A(G5386P1461gat), .B(G5389P1499_bgat), .Y(G5394P1676gat) );
INVXL U_g1730P1422_b (.A(G1730P1422gat), .Y(G1730P1422_bgat) );
OR2XL U_g1899P1680 (.A(G1749P988gat), .B(G1730P1422_bgat), .Y(G1899P1680gat) );
OR2XL U_g1895P1681 (.A(G4716P989gat), .B(G1730P1422_bgat), .Y(G1895P1681gat) );
INVXL U_g1742P992_b (.A(G1742P992gat), .Y(G1742P992_bgat) );
INVXL U_g1856P1513_b (.A(G1856P1513gat), .Y(G1856P1513_bgat) );
AND2XL U_g4708P1684 (.A(G1742P992_bgat), .B(G1856P1513_bgat), .Y(G4708P1684gat) );
OR3XL U_g4700P1685 (.A(G1742P992gat), .B(G1855P1507gat), .C(G1854P1512gat), .Y(G4700P1685gat) );
OR2XL U_g2125P1688 (.A(G1995P993gat), .B(G2124P1506gat), .Y(G2125P1688gat) );
INVXL U_g1064P996_b (.A(G1064P996gat), .Y(G1064P996_bgat) );
INVXL U_g1178P1559_b (.A(G1178P1559gat), .Y(G1178P1559_bgat) );
AND2XL U_g4220P1693 (.A(G1064P996_bgat), .B(G1178P1559_bgat), .Y(G4220P1693gat) );
OR3XL U_g4212P1694 (.A(G1064P996gat), .B(G1177P1524gat), .C(G1176P1558gat), .Y(G4212P1694gat) );
OR2XL U_g1448P1698 (.A(G1318P997gat), .B(G1447P1565gat), .Y(G1448P1698gat) );
INVXL U_g5289P1158_b (.A(G5289P1158gat), .Y(G5289P1158_bgat) );
OR2XL U_g5294P1699 (.A(G5289P1158_bgat), .B(G3350P1331gat), .Y(G5294P1699gat) );
INVXL U_g1301P1000_b (.A(G1301P1000gat), .Y(G1301P1000_bgat) );
INVXL U_g1445P1533_b (.A(G1445P1533gat), .Y(G1445P1533_bgat) );
INVXL U_g1446P1564_b (.A(G1446P1564gat), .Y(G1446P1564_bgat) );
AND3XL U_g4419P1702 (.A(G1301P1000_bgat), .B(G1445P1533_bgat), .C(G1446P1564_bgat), .Y(G4419P1702gat) );
OR4XL U_g4361P1703 (.A(G1301P1000gat), .B(G1444P1531gat), .C(G1442P1535gat), .D(G1443P1562gat), .Y(G4361P1703gat) );
INVXL U_g1046P1001_b (.A(G1046P1001gat), .Y(G1046P1001_bgat) );
INVXL U_g1174P1527_b (.A(G1174P1527gat), .Y(G1174P1527_bgat) );
INVXL U_g1175P1556_b (.A(G1175P1556gat), .Y(G1175P1556_bgat) );
AND3XL U_g4204P1706 (.A(G1046P1001_bgat), .B(G1174P1527_bgat), .C(G1175P1556_bgat), .Y(G4204P1706gat) );
OR4XL U_g4196P1707 (.A(G1046P1001gat), .B(G1173P1523gat), .C(G1171P1526gat), .D(G1172P1557gat), .Y(G4196P1707gat) );
OR5XL U_g1458P1719 (.A(G1341P1010gat), .B(G1456P1578gat), .C(G1455P1585gat), .D(G1454P1593gat), .E(G1457P1597gat), .Y(G1458P1719gat) );
OR5XL U_g1185P1721 (.A(G1097P1011gat), .B(G1183P1568gat), .C(G1182P1588gat), .D(G1181P1590gat), .E(G1184P1604gat), .Y(G1185P1721gat) );
INVXL U_g1052P1426_b (.A(G1052P1426gat), .Y(G1052P1426_bgat) );
OR2XL U_g1221P1722 (.A(G1071P1014gat), .B(G1052P1426_bgat), .Y(G1221P1722gat) );
OR2XL U_g1217P1723 (.A(G4228P1015gat), .B(G1052P1426_bgat), .Y(G1217P1723gat) );
OR3XL U_g4260P1727 (.A(G1145P1020gat), .B(G1195P1605gat), .C(G1196P1651gat), .Y(G4260P1727gat) );
OR2XL U_g1478P1731 (.A(G1404P1021gat), .B(G1477P1600gat), .Y(G1478P1731gat) );
INVXL U_g1382P1024_b (.A(G1382P1024gat), .Y(G1382P1024_bgat) );
INVXL U_g1475P1579_b (.A(G1475P1579gat), .Y(G1475P1579_bgat) );
INVXL U_g1476P1601_b (.A(G1476P1601gat), .Y(G1476P1601_bgat) );
AND3XL U_g4555P1734 (.A(G1382P1024_bgat), .B(G1475P1579_bgat), .C(G1476P1601_bgat), .Y(G4555P1734gat) );
OR4XL U_g4467P1735 (.A(G1382P1024gat), .B(G1474P1573gat), .C(G1472P1580gat), .D(G1473P1599gat), .Y(G4467P1735gat) );
OR4XL U_g4252P1737 (.A(G1128P1025gat), .B(G1192P1569gat), .C(G1193P1606gat), .D(G1194P1652gat), .Y(G4252P1737gat) );
OR5XL U_g4244P1739 (.A(G1111P1028gat), .B(G1189P1567gat), .C(G1188P1587gat), .D(G1190P1603gat), .E(G1191P1649gat), .Y(G4244P1739gat) );
INVXL U_g1359P1029_b (.A(G1359P1029gat), .Y(G1359P1029_bgat) );
INVXL U_g1470P1576_b (.A(G1470P1576gat), .Y(G1470P1576_bgat) );
INVXL U_g1469P1583_b (.A(G1469P1583gat), .Y(G1469P1583_bgat) );
INVXL U_g1471P1598_b (.A(G1471P1598gat), .Y(G1471P1598_bgat) );
AND4XL U_g4575P1742 (.A(G1359P1029_bgat), .B(G1470P1576_bgat), .C(G1469P1583_bgat), .D(G1471P1598_bgat), .Y(G4575P1742gat) );
OR5XL U_g4487P1743 (.A(G1359P1029gat), .B(G1468P1572gat), .C(G1466P1577gat), .D(G1465P1584gat), .E(G1467P1596gat), .Y(G4487P1743gat) );
OR2XL U_g4268P1747 (.A(G1160P1034gat), .B(G1197P1650gat), .Y(G4268P1747gat) );
AND3XL U_g3520P1748 (.A(G3454P1453gat), .B(G3445P1455gat), .C(G3463P1456gat), .Y(G3520P1748gat) );
INVXL U_g3454P1453_b (.A(G3454P1453gat), .Y(G3454P1453_bgat) );
INVXL U_g3445P1455_b (.A(G3445P1455gat), .Y(G3445P1455_bgat) );
AND3XL U_g3523P1749 (.A(G3454P1453_bgat), .B(G3445P1455_bgat), .C(G3463P1456gat), .Y(G3523P1749gat) );
INVXL U_g1812P1404_b (.A(G1812P1404gat), .Y(G1812P1404_bgat) );
OR2XL U_g1929P1751 (.A(G4756P1363gat), .B(G1812P1404_bgat), .Y(G1929P1751gat) );
INVXL U_g5219P1458_b (.A(G5219P1458gat), .Y(G5219P1458_bgat) );
OR2XL U_g5224P1756 (.A(G5219P1458_bgat), .B(G5216P1460gat), .Y(G5224P1756gat) );
INVXL U_g5239P1374_b (.A(G5239P1374gat), .Y(G5239P1374_bgat) );
OR2XL U_g3531P1757 (.A(G5239P1374_bgat), .B(G5236P1457gat), .Y(G3531P1757gat) );
INVXL U_g1852P1149_b (.A(G1852P1149gat), .Y(G1852P1149_bgat) );
INVXL U_g1853P1510_b (.A(G1853P1510gat), .Y(G1853P1510_bgat) );
AND3XL U_g4692P1758 (.A(G3165P927_bgat), .B(G1852P1149_bgat), .C(G1853P1510_bgat), .Y(G4692P1758gat) );
OR4XL U_g4684P1759 (.A(G3165P927gat), .B(G1849P1148gat), .C(G1850P1511gat), .D(G1851P1631gat), .Y(G4684P1759gat) );
INVXL U_g2122P1151_b (.A(G2122P1151gat), .Y(G2122P1151_bgat) );
INVXL U_g2123P1505_b (.A(G2123P1505gat), .Y(G2123P1505_bgat) );
AND3XL U_g4883P1760 (.A(G3165P927_bgat), .B(G2122P1151_bgat), .C(G2123P1505_bgat), .Y(G4883P1760gat) );
OR4XL U_g4825P1761 (.A(G3165P927gat), .B(G2119P1153gat), .C(G2120P1503gat), .D(G2121P1633gat), .Y(G4825P1761gat) );
INVXL U_g5216P1460_b (.A(G5216P1460gat), .Y(G5216P1460_bgat) );
OR2XL U_g5225P1762 (.A(G5219P1458gat), .B(G5216P1460_bgat), .Y(G5225P1762gat) );
AND2XL U_g4111P1765 (.A(G3167P931_bgat), .B(G4107P1644gat), .Y(G4111P1765gat) );
INVXL U_g3468P1469_b (.A(G3468P1469gat), .Y(G3468P1469_bgat) );
INVXL U_g3477P1471_b (.A(G3477P1471gat), .Y(G3477P1471_bgat) );
AND3XL U_g3529P1767 (.A(G3486P1464gat), .B(G3468P1469_bgat), .C(G3477P1471_bgat), .Y(G3529P1767gat) );
INVXL U_g5422P1638_b (.A(G5422P1638gat), .Y(G5422P1638_bgat) );
OR2XL U_g3967P1769 (.A(G5425P1470gat), .B(G5422P1638_bgat), .Y(G3967P1769gat) );
INVXL U_g5229P1467_b (.A(G5229P1467gat), .Y(G5229P1467_bgat) );
OR2XL U_g5234P1771 (.A(G5229P1467_bgat), .B(G5226P1468gat), .Y(G5234P1771gat) );
INVXL U_g5226P1468_b (.A(G5226P1468gat), .Y(G5226P1468_bgat) );
OR2XL U_g5235P1772 (.A(G5229P1467gat), .B(G5226P1468_bgat), .Y(G5235P1772gat) );
AND3XL U_g3526P1773 (.A(G3486P1464gat), .B(G3468P1469gat), .C(G3477P1471gat), .Y(G3526P1773gat) );
AND2XL U_g4112P1774 (.A(G132P60gat), .B(G4107P1644gat), .Y(G4112P1774gat) );
AND2XL U_g1902P1775 (.A(G54P20gat), .B(G1857P1608gat), .Y(G1902P1775gat) );
AND2XL U_g1224P1777 (.A(G4P1gat), .B(G1179P1552gat), .Y(G1224P1777gat) );
INVXL U_g1152P1452_b (.A(G1152P1452gat), .Y(G1152P1452_bgat) );
OR2XL U_g1198P1778 (.A(G4P1gat), .B(G1152P1452_bgat), .Y(G1198P1778gat) );
INVXL U_g4748P1658_b (.A(G4748P1658gat), .Y(G4748P1658_bgat) );
OR2XL U_g1925P1780 (.A(G1794P1406gat), .B(G4748P1658_bgat), .Y(G1925P1780gat) );
INVXL U_g4740P1661_b (.A(G4740P1661gat), .Y(G4740P1661_bgat) );
OR2XL U_g1920P1789 (.A(G1778P1307gat), .B(G4740P1661_bgat), .Y(G1920P1789gat) );
INVXL U_g4732P1670_b (.A(G4732P1670gat), .Y(G4732P1670_bgat) );
OR2XL U_g1915P1790 (.A(G1767P1417gat), .B(G4732P1670_bgat), .Y(G1915P1790gat) );
OR2XL U_g1903P1793 (.A(G1863P1675gat), .B(G1902P1775gat), .Y(G1903P1793gat) );
OR2XL U_g4815P1794 (.A(G2158P1501gat), .B(G2125P1688gat), .Y(G4815P1794gat) );
INVXL U_g1749P988_b (.A(G1749P988gat), .Y(G1749P988_bgat) );
OR2XL U_g1900P1795 (.A(G1749P988_bgat), .B(G1730P1422gat), .Y(G1900P1795gat) );
INVXL U_g4716P989_b (.A(G4716P989gat), .Y(G4716P989_bgat) );
OR2XL U_g1896P1796 (.A(G4716P989_bgat), .B(G1730P1422gat), .Y(G1896P1796gat) );
INVXL U_g4220P1693_b (.A(G4220P1693gat), .Y(G4220P1693_bgat) );
OR2XL U_g1214P1801 (.A(G1034P1429gat), .B(G4220P1693_bgat), .Y(G1214P1801gat) );
INVXL U_g4212P1694_b (.A(G4212P1694gat), .Y(G4212P1694_bgat) );
OR2XL U_g1211P1803 (.A(G1034P1429gat), .B(G4212P1694_bgat), .Y(G1211P1803gat) );
OR2XL U_g4351P1805 (.A(G1481P1528gat), .B(G1448P1698gat), .Y(G4351P1805gat) );
INVXL U_g5295P1536_b (.A(G5295P1536gat), .Y(G5295P1536_bgat) );
INVXL U_g5294P1699_b (.A(G5294P1699gat), .Y(G5294P1699_bgat) );
OR2XL U_g5376P1808 (.A(G5295P1536_bgat), .B(G5294P1699_bgat), .Y(G5376P1808gat) );
INVXL U_g4204P1706_b (.A(G4204P1706gat), .Y(G4204P1706_bgat) );
OR2XL U_g1207P1811 (.A(G1023P1432gat), .B(G4204P1706_bgat), .Y(G1207P1811gat) );
INVXL U_g4196P1707_b (.A(G4196P1707gat), .Y(G4196P1707_bgat) );
OR2XL U_g1204P1813 (.A(G1023P1432gat), .B(G4196P1707_bgat), .Y(G1204P1813gat) );
INVXL U_g4244P1739_b (.A(G4244P1739gat), .Y(G4244P1739_bgat) );
OR2XL U_g1237P1818 (.A(G1089P1436gat), .B(G4244P1739_bgat), .Y(G1237P1818gat) );
OR2XL U_g1225P1819 (.A(G1185P1721gat), .B(G1224P1777gat), .Y(G1225P1819gat) );
INVXL U_g1071P1014_b (.A(G1071P1014gat), .Y(G1071P1014_bgat) );
OR2XL U_g1222P1820 (.A(G1071P1014_bgat), .B(G1052P1426gat), .Y(G1222P1820gat) );
INVXL U_g4228P1015_b (.A(G4228P1015gat), .Y(G4228P1015_bgat) );
OR2XL U_g1218P1821 (.A(G4228P1015_bgat), .B(G1052P1426gat), .Y(G1218P1821gat) );
INVXL U_g4260P1727_b (.A(G4260P1727gat), .Y(G4260P1727_bgat) );
OR2XL U_g1247P1822 (.A(G1116P1446gat), .B(G4260P1727_bgat), .Y(G1247P1822gat) );
INVXL U_g4268P1747_b (.A(G4268P1747gat), .Y(G4268P1747_bgat) );
OR2XL U_g1252P1824 (.A(G1134P1442gat), .B(G4268P1747_bgat), .Y(G1252P1824gat) );
OR2XL U_g4477P1825 (.A(G1482P1575gat), .B(G1478P1731gat), .Y(G4477P1825gat) );
INVXL U_g4252P1737_b (.A(G4252P1737gat), .Y(G4252P1737_bgat) );
OR2XL U_g1242P1829 (.A(G1100P1448gat), .B(G4252P1737_bgat), .Y(G1242P1829gat) );
INVXL U_g3852P1190_b (.A(G3852P1190gat), .Y(G3852P1190_bgat) );
AND3XL U_g3943P1834 (.A(G3852P1190_bgat), .B(G3871P1548gat), .C(G3862P1566gat), .Y(G3943P1834gat) );
INVXL U_g3862P1566_b (.A(G3862P1566gat), .Y(G3862P1566_bgat) );
AND3XL U_g3946P1835 (.A(G3852P1190gat), .B(G3871P1548gat), .C(G3862P1566_bgat), .Y(G3946P1835gat) );
INVXL U_g4467P1735_b (.A(G4467P1735gat), .Y(G4467P1735_bgat) );
OR2XL U_g4472P1836 (.A(G4464P1032gat), .B(G4467P1735_bgat), .Y(G4472P1836gat) );
INVXL U_g4555P1734_b (.A(G4555P1734gat), .Y(G4555P1734_bgat) );
OR2XL U_g4560P1837 (.A(G1412P1033gat), .B(G4555P1734_bgat), .Y(G4560P1837gat) );
INVXL U_g3463P1456_b (.A(G3463P1456gat), .Y(G3463P1456_bgat) );
AND3XL U_g3519P1839 (.A(G3454P1453gat), .B(G3445P1455_bgat), .C(G3463P1456_bgat), .Y(G3519P1839gat) );
INVXL U_g4756P1363_b (.A(G4756P1363gat), .Y(G4756P1363_bgat) );
OR2XL U_g1930P1840 (.A(G4756P1363_bgat), .B(G1812P1404gat), .Y(G1930P1840gat) );
INVXL U_g5009P1664_b (.A(G5009P1664gat), .Y(G5009P1664_bgat) );
OR2XL U_g5014P1841 (.A(G3137P914gat), .B(G5009P1664_bgat), .Y(G5014P1841gat) );
OR2XL U_g4931P1842 (.A(G2159P1621gat), .B(G2155P1657gat), .Y(G4931P1842gat) );
AND3XL U_g3949P1843 (.A(G3328P916gat), .B(G3883P1473gat), .C(G3892P1490gat), .Y(G3949P1843gat) );
INVXL U_g3328P916_b (.A(G3328P916gat), .Y(G3328P916_bgat) );
INVXL U_g3883P1473_b (.A(G3883P1473gat), .Y(G3883P1473_bgat) );
AND3XL U_g3952P1844 (.A(G3328P916_bgat), .B(G3883P1473_bgat), .C(G3892P1490gat), .Y(G3952P1844gat) );
AND3XL U_g3522P1845 (.A(G3454P1453_bgat), .B(G3445P1455gat), .C(G3463P1456_bgat), .Y(G3522P1845gat) );
INVXL U_g5224P1756_b (.A(G5224P1756gat), .Y(G5224P1756_bgat) );
INVXL U_g5225P1762_b (.A(G5225P1762gat), .Y(G5225P1762_bgat) );
OR2XL U_g5247P1847 (.A(G5224P1756_bgat), .B(G5225P1762_bgat), .Y(G5247P1847gat) );
INVXL U_g4708P1684_b (.A(G4708P1684gat), .Y(G4708P1684_bgat) );
OR2XL U_g1892P1848 (.A(G3165P927_bgat), .B(G4708P1684_bgat), .Y(G1892P1848gat) );
INVXL U_g4700P1685_b (.A(G4700P1685gat), .Y(G4700P1685_bgat) );
OR2XL U_g1889P1850 (.A(G3165P927_bgat), .B(G4700P1685_bgat), .Y(G1889P1850gat) );
INVXL U_g5386P1461_b (.A(G5386P1461gat), .Y(G5386P1461_bgat) );
OR2XL U_g5395P1856 (.A(G5386P1461_bgat), .B(G5389P1499gat), .Y(G5395P1856gat) );
INVXL U_g4684P1759_b (.A(G4684P1759gat), .Y(G4684P1759_bgat) );
OR2XL U_g1882P1857 (.A(G3167P931_bgat), .B(G4684P1759_bgat), .Y(G1882P1857gat) );
INVXL U_g4692P1758_b (.A(G4692P1758gat), .Y(G4692P1758_bgat) );
OR2XL U_g1885P1858 (.A(G3167P931_bgat), .B(G4692P1758_bgat), .Y(G1885P1858gat) );
OR2XL U_g4113P1859 (.A(G4111P1765gat), .B(G4112P1774gat), .Y(G4113P1859gat) );
INVXL U_g5234P1771_b (.A(G5234P1771gat), .Y(G5234P1771_bgat) );
INVXL U_g5235P1772_b (.A(G5235P1772gat), .Y(G5235P1772_bgat) );
OR2XL U_g5255P1860 (.A(G5234P1771_bgat), .B(G5235P1772_bgat), .Y(G5255P1860gat) );
INVXL U_g3486P1464_b (.A(G3486P1464gat), .Y(G3486P1464_bgat) );
AND3XL U_g3528P1861 (.A(G3486P1464_bgat), .B(G3468P1469gat), .C(G3477P1471_bgat), .Y(G3528P1861gat) );
INVXL U_g5425P1470_b (.A(G5425P1470gat), .Y(G5425P1470_bgat) );
OR2XL U_g3966P1862 (.A(G5425P1470_bgat), .B(G5422P1638gat), .Y(G3966P1862gat) );
AND3XL U_g3525P1863 (.A(G3486P1464_bgat), .B(G3468P1469_bgat), .C(G3477P1471gat), .Y(G3525P1863gat) );
INVXL U_g4P1_b (.A(G4P1gat), .Y(G4P1_bgat) );
OR2XL U_g1199P1865 (.A(G4P1_bgat), .B(G1152P1452gat), .Y(G1199P1865gat) );
AND3XL U_g3733P1868 (.A(G3717P169_bgat), .B(G3724P170gat), .C(G4113P1859gat), .Y(G3733P1868gat) );
INVXL U_g1694P160_b (.A(G1694P160gat), .Y(G1694P160_bgat) );
AND3XL U_g2335P1869 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G3848P1864gat), .Y(G2335P1869gat) );
INVXL U_g1690P158_b (.A(G1690P158gat), .Y(G1690P158_bgat) );
AND3XL U_g1664P1870 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G3848P1864gat), .Y(G1664P1870gat) );
INVXL U_g1794P1406_b (.A(G1794P1406gat), .Y(G1794P1406_bgat) );
OR2XL U_g1924P1872 (.A(G1794P1406_bgat), .B(G4748P1658gat), .Y(G1924P1872gat) );
INVXL U_g4931P1842_b (.A(G4931P1842gat), .Y(G4931P1842_bgat) );
OR2XL U_g4936P1873 (.A(G4928P1665gat), .B(G4931P1842_bgat), .Y(G4936P1873gat) );
INVXL U_g1778P1307_b (.A(G1778P1307gat), .Y(G1778P1307_bgat) );
OR2XL U_g1919P1874 (.A(G1778P1307_bgat), .B(G4740P1661gat), .Y(G1919P1874gat) );
INVXL U_g1767P1417_b (.A(G1767P1417gat), .Y(G1767P1417_bgat) );
OR2XL U_g1914P1875 (.A(G1767P1417_bgat), .B(G4732P1670gat), .Y(G1914P1875gat) );
INVXL U_g5394P1676_b (.A(G5394P1676gat), .Y(G5394P1676_bgat) );
INVXL U_g5395P1856_b (.A(G5395P1856gat), .Y(G5395P1856_bgat) );
OR2XL U_g5417P1877 (.A(G5394P1676_bgat), .B(G5395P1856_bgat), .Y(G5417P1877gat) );
INVXL U_g4815P1794_b (.A(G4815P1794gat), .Y(G4815P1794_bgat) );
OR2XL U_g4820P1879 (.A(G4812P986gat), .B(G4815P1794_bgat), .Y(G4820P1879gat) );
OR2XL U_g4878P1880 (.A(G2001P987gat), .B(G2125P1688gat), .Y(G4878P1880gat) );
INVXL U_g1758P1420_b (.A(G1758P1420gat), .Y(G1758P1420_bgat) );
AND2XL U_g1953P1881 (.A(G1758P1420_bgat), .B(G1903P1793gat), .Y(G1953P1881gat) );
INVXL U_g1899P1680_b (.A(G1899P1680gat), .Y(G1899P1680_bgat) );
INVXL U_g1900P1795_b (.A(G1900P1795gat), .Y(G1900P1795_bgat) );
OR2XL U_g1901P1882 (.A(G1899P1680_bgat), .B(G1900P1795_bgat), .Y(G1901P1882gat) );
INVXL U_g1895P1681_b (.A(G1895P1681gat), .Y(G1895P1681_bgat) );
INVXL U_g1896P1796_b (.A(G1896P1796gat), .Y(G1896P1796_bgat) );
OR2XL U_g1897P1883 (.A(G1895P1681_bgat), .B(G1896P1796_bgat), .Y(G1897P1883gat) );
INVXL U_g5376P1808_b (.A(G5376P1808gat), .Y(G5376P1808_bgat) );
OR2XL U_g5385P1885 (.A(G5379P1518gat), .B(G5376P1808_bgat), .Y(G5385P1885gat) );
INVXL U_g1034P1429_b (.A(G1034P1429gat), .Y(G1034P1429_bgat) );
OR2XL U_g1213P1889 (.A(G1034P1429_bgat), .B(G4220P1693gat), .Y(G1213P1889gat) );
OR2XL U_g1210P1890 (.A(G1034P1429_bgat), .B(G4212P1694gat), .Y(G1210P1890gat) );
INVXL U_g1023P1432_b (.A(G1023P1432gat), .Y(G1023P1432_bgat) );
OR2XL U_g1203P1891 (.A(G1023P1432_bgat), .B(G4196P1707gat), .Y(G1203P1891gat) );
OR2XL U_g1206P1892 (.A(G1023P1432_bgat), .B(G4204P1706gat), .Y(G1206P1892gat) );
INVXL U_g1451P1551_b (.A(G1451P1551gat), .Y(G1451P1551_bgat) );
INVXL U_g1458P1719_b (.A(G1458P1719gat), .Y(G1458P1719_bgat) );
AND2XL U_g1483P1895 (.A(G1451P1551_bgat), .B(G1458P1719_bgat), .Y(G1483P1895gat) );
INVXL U_g1089P1436_b (.A(G1089P1436gat), .Y(G1089P1436_bgat) );
OR2XL U_g1236P1896 (.A(G1089P1436_bgat), .B(G4244P1739gat), .Y(G1236P1896gat) );
INVXL U_g1080P1438_b (.A(G1080P1438gat), .Y(G1080P1438_bgat) );
AND2XL U_g1272P1898 (.A(G1080P1438_bgat), .B(G1225P1819gat), .Y(G1272P1898gat) );
INVXL U_g1221P1722_b (.A(G1221P1722gat), .Y(G1221P1722_bgat) );
INVXL U_g1222P1820_b (.A(G1222P1820gat), .Y(G1222P1820_bgat) );
OR2XL U_g1223P1899 (.A(G1221P1722_bgat), .B(G1222P1820_bgat), .Y(G1223P1899gat) );
INVXL U_g1217P1723_b (.A(G1217P1723gat), .Y(G1217P1723_bgat) );
INVXL U_g1218P1821_b (.A(G1218P1821gat), .Y(G1218P1821_bgat) );
OR2XL U_g1219P1900 (.A(G1217P1723_bgat), .B(G1218P1821_bgat), .Y(G1219P1900gat) );
INVXL U_g4351P1805_b (.A(G4351P1805gat), .Y(G4351P1805_bgat) );
OR2XL U_g4356P1901 (.A(G4348P1016gat), .B(G4351P1805_bgat), .Y(G4356P1901gat) );
OR2XL U_g4414P1902 (.A(G1324P1017gat), .B(G1448P1698gat), .Y(G4414P1902gat) );
INVXL U_g1134P1442_b (.A(G1134P1442gat), .Y(G1134P1442_bgat) );
OR2XL U_g1251P1903 (.A(G1134P1442_bgat), .B(G4268P1747gat), .Y(G1251P1903gat) );
INVXL U_g1116P1446_b (.A(G1116P1446gat), .Y(G1116P1446_bgat) );
OR2XL U_g1246P1906 (.A(G1116P1446_bgat), .B(G4260P1727gat), .Y(G1246P1906gat) );
INVXL U_g1100P1448_b (.A(G1100P1448gat), .Y(G1100P1448_bgat) );
OR2XL U_g1241P1907 (.A(G1100P1448_bgat), .B(G4252P1737gat), .Y(G1241P1907gat) );
INVXL U_g3871P1548_b (.A(G3871P1548gat), .Y(G3871P1548_bgat) );
AND3XL U_g3945P1908 (.A(G3852P1190_bgat), .B(G3871P1548_bgat), .C(G3862P1566_bgat), .Y(G3945P1908gat) );
AND3XL U_g3942P1909 (.A(G3852P1190gat), .B(G3871P1548_bgat), .C(G3862P1566gat), .Y(G3942P1909gat) );
INVXL U_g4464P1032_b (.A(G4464P1032gat), .Y(G4464P1032_bgat) );
OR2XL U_g4473P1910 (.A(G4464P1032_bgat), .B(G4467P1735gat), .Y(G4473P1910gat) );
INVXL U_g1412P1033_b (.A(G1412P1033gat), .Y(G1412P1033_bgat) );
OR2XL U_g4561P1911 (.A(G1412P1033_bgat), .B(G4555P1734gat), .Y(G4561P1911gat) );
INVXL U_g3520P1748_b (.A(G3520P1748gat), .Y(G3520P1748_bgat) );
INVXL U_g3519P1839_b (.A(G3519P1839gat), .Y(G3519P1839_bgat) );
AND2XL U_g3521P1912 (.A(G3520P1748_bgat), .B(G3519P1839_bgat), .Y(G3521P1912gat) );
INVXL U_g3523P1749_b (.A(G3523P1749gat), .Y(G3523P1749_bgat) );
INVXL U_g3522P1845_b (.A(G3522P1845gat), .Y(G3522P1845_bgat) );
AND2XL U_g3524P1913 (.A(G3523P1749_bgat), .B(G3522P1845_bgat), .Y(G3524P1913gat) );
INVXL U_g1929P1751_b (.A(G1929P1751gat), .Y(G1929P1751_bgat) );
INVXL U_g1930P1840_b (.A(G1930P1840gat), .Y(G1930P1840_bgat) );
OR2XL U_g1931P1914 (.A(G1929P1751_bgat), .B(G1930P1840_bgat), .Y(G1931P1914gat) );
OR2XL U_g5015P1915 (.A(G3137P914_bgat), .B(G5009P1664gat), .Y(G5015P1915gat) );
INVXL U_g2128P1619_b (.A(G2128P1619gat), .Y(G2128P1619_bgat) );
INVXL U_g2135P1673_b (.A(G2135P1673gat), .Y(G2135P1673_bgat) );
AND2XL U_g2160P1916 (.A(G2128P1619_bgat), .B(G2135P1673_bgat), .Y(G2160P1916gat) );
INVXL U_g3892P1490_b (.A(G3892P1490gat), .Y(G3892P1490_bgat) );
AND3XL U_g3951P1918 (.A(G3328P916gat), .B(G3883P1473_bgat), .C(G3892P1490_bgat), .Y(G3951P1918gat) );
AND3XL U_g3948P1919 (.A(G3328P916_bgat), .B(G3883P1473gat), .C(G3892P1490_bgat), .Y(G3948P1919gat) );
OR2XL U_g1891P1923 (.A(G3165P927gat), .B(G4708P1684gat), .Y(G1891P1923gat) );
OR2XL U_g1888P1924 (.A(G3165P927gat), .B(G4700P1685gat), .Y(G1888P1924gat) );
OR2XL U_g1881P1927 (.A(G3167P931gat), .B(G4684P1759gat), .Y(G1881P1927gat) );
OR2XL U_g1884P1928 (.A(G3167P931gat), .B(G4692P1758gat), .Y(G1884P1928gat) );
INVXL U_g3529P1767_b (.A(G3529P1767gat), .Y(G3529P1767_bgat) );
INVXL U_g3528P1861_b (.A(G3528P1861gat), .Y(G3528P1861_bgat) );
AND2XL U_g3530P1929 (.A(G3529P1767_bgat), .B(G3528P1861_bgat), .Y(G3530P1929gat) );
INVXL U_g3526P1773_b (.A(G3526P1773gat), .Y(G3526P1773_bgat) );
INVXL U_g3525P1863_b (.A(G3525P1863gat), .Y(G3525P1863_bgat) );
AND2XL U_g3527P1932 (.A(G3526P1773_bgat), .B(G3525P1863_bgat), .Y(G3527P1932gat) );
INVXL U_g1198P1778_b (.A(G1198P1778gat), .Y(G1198P1778_bgat) );
INVXL U_g1199P1865_b (.A(G1199P1865gat), .Y(G1199P1865_bgat) );
OR2XL U_g1200P1934 (.A(G1198P1778_bgat), .B(G1199P1865_bgat), .Y(G1200P1934gat) );
AND3XL U_g3840P1935 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1931P1914gat), .Y(G3840P1935gat) );
AND3XL U_g3779P1936 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1200P1934gat), .Y(G3779P1936gat) );
INVXL U_g1925P1780_b (.A(G1925P1780gat), .Y(G1925P1780_bgat) );
INVXL U_g1924P1872_b (.A(G1924P1872gat), .Y(G1924P1872_bgat) );
OR2XL U_g1926P1937 (.A(G1925P1780_bgat), .B(G1924P1872_bgat), .Y(G1926P1937gat) );
INVXL U_g4928P1665_b (.A(G4928P1665gat), .Y(G4928P1665_bgat) );
OR2XL U_g4937P1938 (.A(G4928P1665_bgat), .B(G4931P1842gat), .Y(G4937P1938gat) );
INVXL U_g1920P1789_b (.A(G1920P1789gat), .Y(G1920P1789_bgat) );
INVXL U_g1919P1874_b (.A(G1919P1874gat), .Y(G1919P1874_bgat) );
OR2XL U_g1921P1939 (.A(G1920P1789_bgat), .B(G1919P1874_bgat), .Y(G1921P1939gat) );
INVXL U_g1915P1790_b (.A(G1915P1790gat), .Y(G1915P1790_bgat) );
INVXL U_g1914P1875_b (.A(G1914P1875gat), .Y(G1914P1875_bgat) );
OR2XL U_g1916P1940 (.A(G1915P1790_bgat), .B(G1914P1875_bgat), .Y(G1916P1940gat) );
INVXL U_g1903P1793_b (.A(G1903P1793gat), .Y(G1903P1793_bgat) );
AND2XL U_g1947P1941 (.A(G1903P1793_bgat), .B(G1901P1882gat), .Y(G1947P1941gat) );
INVXL U_g4812P986_b (.A(G4812P986gat), .Y(G4812P986_bgat) );
OR2XL U_g4821P1943 (.A(G4812P986_bgat), .B(G4815P1794gat), .Y(G4821P1943gat) );
INVXL U_g2001P987_b (.A(G2001P987gat), .Y(G2001P987_bgat) );
INVXL U_g2125P1688_b (.A(G2125P1688gat), .Y(G2125P1688_bgat) );
OR2XL U_g4879P1944 (.A(G2001P987_bgat), .B(G2125P1688_bgat), .Y(G4879P1944gat) );
AND2XL U_g1952P1945 (.A(G1758P1420gat), .B(G1903P1793_bgat), .Y(G1952P1945gat) );
INVXL U_g5379P1518_b (.A(G5379P1518gat), .Y(G5379P1518_bgat) );
OR2XL U_g5384P1947 (.A(G5379P1518_bgat), .B(G5376P1808gat), .Y(G5384P1947gat) );
INVXL U_g1214P1801_b (.A(G1214P1801gat), .Y(G1214P1801_bgat) );
INVXL U_g1213P1889_b (.A(G1213P1889gat), .Y(G1213P1889_bgat) );
OR2XL U_g1215P1948 (.A(G1214P1801_bgat), .B(G1213P1889_bgat), .Y(G1215P1948gat) );
INVXL U_g1211P1803_b (.A(G1211P1803gat), .Y(G1211P1803_bgat) );
INVXL U_g1210P1890_b (.A(G1210P1890gat), .Y(G1210P1890_bgat) );
OR2XL U_g1212P1949 (.A(G1211P1803_bgat), .B(G1210P1890_bgat), .Y(G1212P1949gat) );
INVXL U_g1207P1811_b (.A(G1207P1811gat), .Y(G1207P1811_bgat) );
INVXL U_g1206P1892_b (.A(G1206P1892gat), .Y(G1206P1892_bgat) );
OR2XL U_g1208P1950 (.A(G1207P1811_bgat), .B(G1206P1892_bgat), .Y(G1208P1950gat) );
INVXL U_g1204P1813_b (.A(G1204P1813gat), .Y(G1204P1813_bgat) );
INVXL U_g1203P1891_b (.A(G1203P1891gat), .Y(G1203P1891_bgat) );
OR2XL U_g1205P1951 (.A(G1204P1813_bgat), .B(G1203P1891_bgat), .Y(G1205P1951gat) );
INVXL U_g1237P1818_b (.A(G1237P1818gat), .Y(G1237P1818_bgat) );
INVXL U_g1236P1896_b (.A(G1236P1896gat), .Y(G1236P1896_bgat) );
OR2XL U_g1238P1953 (.A(G1237P1818_bgat), .B(G1236P1896_bgat), .Y(G1238P1953gat) );
INVXL U_g1225P1819_b (.A(G1225P1819gat), .Y(G1225P1819_bgat) );
AND2XL U_g1266P1954 (.A(G1225P1819_bgat), .B(G1223P1899gat), .Y(G1266P1954gat) );
AND2XL U_g1271P1955 (.A(G1080P1438gat), .B(G1225P1819_bgat), .Y(G1271P1955gat) );
INVXL U_g4348P1016_b (.A(G4348P1016gat), .Y(G4348P1016_bgat) );
OR2XL U_g4357P1957 (.A(G4348P1016_bgat), .B(G4351P1805gat), .Y(G4357P1957gat) );
INVXL U_g1324P1017_b (.A(G1324P1017gat), .Y(G1324P1017_bgat) );
INVXL U_g1448P1698_b (.A(G1448P1698gat), .Y(G1448P1698_bgat) );
OR2XL U_g4415P1958 (.A(G1324P1017_bgat), .B(G1448P1698_bgat), .Y(G4415P1958gat) );
INVXL U_g1247P1822_b (.A(G1247P1822gat), .Y(G1247P1822_bgat) );
INVXL U_g1246P1906_b (.A(G1246P1906gat), .Y(G1246P1906_bgat) );
OR2XL U_g1248P1959 (.A(G1247P1822_bgat), .B(G1246P1906_bgat), .Y(G1248P1959gat) );
INVXL U_g1252P1824_b (.A(G1252P1824gat), .Y(G1252P1824_bgat) );
INVXL U_g1251P1903_b (.A(G1251P1903gat), .Y(G1251P1903_bgat) );
OR2XL U_g1253P1960 (.A(G1252P1824_bgat), .B(G1251P1903_bgat), .Y(G1253P1960gat) );
INVXL U_g1242P1829_b (.A(G1242P1829gat), .Y(G1242P1829_bgat) );
INVXL U_g1241P1907_b (.A(G1241P1907gat), .Y(G1241P1907_bgat) );
OR2XL U_g1243P1961 (.A(G1242P1829_bgat), .B(G1241P1907_bgat), .Y(G1243P1961gat) );
INVXL U_g3943P1834_b (.A(G3943P1834gat), .Y(G3943P1834_bgat) );
INVXL U_g3942P1909_b (.A(G3942P1909gat), .Y(G3942P1909_bgat) );
AND2XL U_g3944P1962 (.A(G3943P1834_bgat), .B(G3942P1909_bgat), .Y(G3944P1962gat) );
INVXL U_g3946P1835_b (.A(G3946P1835gat), .Y(G3946P1835_bgat) );
INVXL U_g3945P1908_b (.A(G3945P1908gat), .Y(G3945P1908_bgat) );
AND2XL U_g3947P1963 (.A(G3946P1835_bgat), .B(G3945P1908_bgat), .Y(G3947P1963gat) );
INVXL U_g4472P1836_b (.A(G4472P1836gat), .Y(G4472P1836_bgat) );
INVXL U_g4473P1910_b (.A(G4473P1910gat), .Y(G4473P1910_bgat) );
OR2XL U_g4474P1964 (.A(G4472P1836_bgat), .B(G4473P1910_bgat), .Y(G4474P1964gat) );
INVXL U_g4560P1837_b (.A(G4560P1837gat), .Y(G4560P1837_bgat) );
INVXL U_g4561P1911_b (.A(G4561P1911gat), .Y(G4561P1911_bgat) );
OR2XL U_g4562P1965 (.A(G4560P1837_bgat), .B(G4561P1911_bgat), .Y(G4562P1965gat) );
INVXL U_g3521P1912_b (.A(G3521P1912gat), .Y(G3521P1912_bgat) );
INVXL U_g3524P1913_b (.A(G3524P1913gat), .Y(G3524P1913_bgat) );
OR2XL U_g5244P1966 (.A(G3521P1912_bgat), .B(G3524P1913_bgat), .Y(G5244P1966gat) );
INVXL U_g5014P1841_b (.A(G5014P1841gat), .Y(G5014P1841_bgat) );
INVXL U_g5015P1915_b (.A(G5015P1915gat), .Y(G5015P1915_bgat) );
OR2XL U_g5016P1968 (.A(G5014P1841_bgat), .B(G5015P1915_bgat), .Y(G5016P1968gat) );
INVXL U_g3949P1843_b (.A(G3949P1843gat), .Y(G3949P1843_bgat) );
INVXL U_g3948P1919_b (.A(G3948P1919gat), .Y(G3948P1919_bgat) );
AND2XL U_g3950P1970 (.A(G3949P1843_bgat), .B(G3948P1919_bgat), .Y(G3950P1970gat) );
INVXL U_g3952P1844_b (.A(G3952P1844gat), .Y(G3952P1844_bgat) );
INVXL U_g3951P1918_b (.A(G3951P1918gat), .Y(G3951P1918_bgat) );
AND2XL U_g3953P1971 (.A(G3952P1844_bgat), .B(G3951P1918_bgat), .Y(G3953P1971gat) );
INVXL U_g1892P1848_b (.A(G1892P1848gat), .Y(G1892P1848_bgat) );
INVXL U_g1891P1923_b (.A(G1891P1923gat), .Y(G1891P1923_bgat) );
OR2XL U_g1893P1972 (.A(G1892P1848_bgat), .B(G1891P1923_bgat), .Y(G1893P1972gat) );
INVXL U_g1889P1850_b (.A(G1889P1850gat), .Y(G1889P1850_bgat) );
INVXL U_g1888P1924_b (.A(G1888P1924gat), .Y(G1888P1924_bgat) );
OR2XL U_g1890P1973 (.A(G1889P1850_bgat), .B(G1888P1924_bgat), .Y(G1890P1973gat) );
INVXL U_g1882P1857_b (.A(G1882P1857gat), .Y(G1882P1857_bgat) );
INVXL U_g1881P1927_b (.A(G1881P1927gat), .Y(G1881P1927_bgat) );
OR2XL U_g1883P1974 (.A(G1882P1857_bgat), .B(G1881P1927_bgat), .Y(G1883P1974gat) );
INVXL U_g1885P1858_b (.A(G1885P1858gat), .Y(G1885P1858_bgat) );
INVXL U_g1884P1928_b (.A(G1884P1928gat), .Y(G1884P1928_bgat) );
OR2XL U_g1886P1975 (.A(G1885P1858_bgat), .B(G1884P1928_bgat), .Y(G1886P1975gat) );
INVXL U_g3530P1929_b (.A(G3530P1929gat), .Y(G3530P1929_bgat) );
INVXL U_g3527P1932_b (.A(G3527P1932gat), .Y(G3527P1932_bgat) );
OR2XL U_g5252P1976 (.A(G3530P1929_bgat), .B(G3527P1932_bgat), .Y(G5252P1976gat) );
AND3XL U_g4068P1980 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1916P1940gat), .Y(G4068P1980gat) );
AND3XL U_g4010P1981 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1238P1953gat), .Y(G4010P1981gat) );
AND3XL U_g3846P1982 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1921P1939gat), .Y(G3846P1982gat) );
AND3XL U_g3843P1983 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1926P1937gat), .Y(G3843P1983gat) );
AND3XL U_g3788P1984 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1243P1961gat), .Y(G3788P1984gat) );
AND3XL U_g3785P1985 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1248P1959gat), .Y(G3785P1985gat) );
AND3XL U_g3782P1986 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1253P1960gat), .Y(G3782P1986gat) );
INVXL U_g2155P1657_b (.A(G2155P1657gat), .Y(G2155P1657_bgat) );
INVXL U_g5016P1968_b (.A(G5016P1968gat), .Y(G5016P1968_bgat) );
OR2XL U_g5025P1987 (.A(G2155P1657_bgat), .B(G5016P1968_bgat), .Y(G5025P1987gat) );
INVXL U_g4936P1873_b (.A(G4936P1873gat), .Y(G4936P1873_bgat) );
INVXL U_g4937P1938_b (.A(G4937P1938gat), .Y(G4937P1938_bgat) );
OR2XL U_g4938P1989 (.A(G4936P1873_bgat), .B(G4937P1938_bgat), .Y(G4938P1989gat) );
AND2XL U_g1943P1992 (.A(G1903P1793gat), .B(G1890P1973gat), .Y(G1943P1992gat) );
INVXL U_g1897P1883_b (.A(G1897P1883gat), .Y(G1897P1883_bgat) );
AND2XL U_g1948P1993 (.A(G1903P1793gat), .B(G1897P1883_bgat), .Y(G1948P1993gat) );
AND2XL U_g1935P1994 (.A(G1903P1793gat), .B(G1883P1974gat), .Y(G1935P1994gat) );
INVXL U_g4820P1879_b (.A(G4820P1879gat), .Y(G4820P1879_bgat) );
INVXL U_g4821P1943_b (.A(G4821P1943gat), .Y(G4821P1943_bgat) );
OR2XL U_g4822P1995 (.A(G4820P1879_bgat), .B(G4821P1943_bgat), .Y(G4822P1995gat) );
INVXL U_g4878P1880_b (.A(G4878P1880gat), .Y(G4878P1880_bgat) );
INVXL U_g4879P1944_b (.A(G4879P1944gat), .Y(G4879P1944_bgat) );
OR2XL U_g4880P1996 (.A(G4878P1880_bgat), .B(G4879P1944_bgat), .Y(G4880P1996gat) );
OR2XL U_g1954P1997 (.A(G1953P1881gat), .B(G1952P1945gat), .Y(G1954P1997gat) );
INVXL U_g5385P1885_b (.A(G5385P1885gat), .Y(G5385P1885_bgat) );
INVXL U_g5384P1947_b (.A(G5384P1947gat), .Y(G5384P1947_bgat) );
OR2XL U_g5409P1998 (.A(G5385P1885_bgat), .B(G5384P1947_bgat), .Y(G5409P1998gat) );
AND2XL U_g1262P2002 (.A(G1225P1819gat), .B(G1212P1949gat), .Y(G1262P2002gat) );
INVXL U_g1219P1900_b (.A(G1219P1900gat), .Y(G1219P1900_bgat) );
AND2XL U_g1267P2003 (.A(G1225P1819gat), .B(G1219P1900_bgat), .Y(G1267P2003gat) );
AND2XL U_g1257P2004 (.A(G1225P1819gat), .B(G1205P1951gat), .Y(G1257P2004gat) );
OR2XL U_g1273P2005 (.A(G1272P1898gat), .B(G1271P1955gat), .Y(G1273P2005gat) );
INVXL U_g4356P1901_b (.A(G4356P1901gat), .Y(G4356P1901_bgat) );
INVXL U_g4357P1957_b (.A(G4357P1957gat), .Y(G4357P1957_bgat) );
OR2XL U_g4358P2006 (.A(G4356P1901_bgat), .B(G4357P1957_bgat), .Y(G4358P2006gat) );
INVXL U_g4414P1902_b (.A(G4414P1902gat), .Y(G4414P1902_bgat) );
INVXL U_g4415P1958_b (.A(G4415P1958gat), .Y(G4415P1958_bgat) );
OR2XL U_g4416P2007 (.A(G4414P1902_bgat), .B(G4415P1958_bgat), .Y(G4416P2007gat) );
INVXL U_g4474P1964_b (.A(G4474P1964gat), .Y(G4474P1964_bgat) );
OR2XL U_g4483P2010 (.A(G4477P1825gat), .B(G4474P1964_bgat), .Y(G4483P2010gat) );
INVXL U_g1478P1731_b (.A(G1478P1731gat), .Y(G1478P1731_bgat) );
INVXL U_g4562P1965_b (.A(G4562P1965gat), .Y(G4562P1965_bgat) );
OR2XL U_g4571P2011 (.A(G1478P1731_bgat), .B(G4562P1965_bgat), .Y(G4571P2011gat) );
INVXL U_g3944P1962_b (.A(G3944P1962gat), .Y(G3944P1962_bgat) );
INVXL U_g3947P1963_b (.A(G3947P1963gat), .Y(G3947P1963_bgat) );
OR2XL U_g5406P2013 (.A(G3944P1962_bgat), .B(G3947P1963_bgat), .Y(G5406P2013gat) );
INVXL U_g3950P1970_b (.A(G3950P1970gat), .Y(G3950P1970_bgat) );
INVXL U_g3953P1971_b (.A(G3953P1971gat), .Y(G3953P1971_bgat) );
OR2XL U_g5414P2018 (.A(G3950P1970_bgat), .B(G3953P1971_bgat), .Y(G5414P2018gat) );
INVXL U_g5244P1966_b (.A(G5244P1966gat), .Y(G5244P1966_bgat) );
OR2XL U_g3537P2019 (.A(G5247P1847gat), .B(G5244P1966_bgat), .Y(G3537P2019gat) );
INVXL U_g5252P1976_b (.A(G5252P1976gat), .Y(G5252P1976_bgat) );
OR2XL U_g3542P2023 (.A(G5255P1860gat), .B(G5252P1976_bgat), .Y(G3542P2023gat) );
AND3XL U_g4071P2026 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1954P1997gat), .Y(G4071P2026gat) );
AND3XL U_g4013P2027 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1273P2005gat), .Y(G4013P2027gat) );
AND3XL U_g2341P2032 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G3849P2024gat), .Y(G2341P2032gat) );
AND3XL U_g2337P2033 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G3790P2025gat), .Y(G2337P2033gat) );
AND3XL U_g1670P2034 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G3849P2024gat), .Y(G1670P2034gat) );
AND3XL U_g1666P2035 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G3790P2025gat), .Y(G1666P2035gat) );
OR2XL U_g5024P2036 (.A(G2155P1657gat), .B(G5016P1968gat), .Y(G5024P2036gat) );
INVXL U_g4938P1989_b (.A(G4938P1989gat), .Y(G4938P1989_bgat) );
OR2XL U_g4947P2038 (.A(G4941P1669gat), .B(G4938P1989_bgat), .Y(G4947P2038gat) );
INVXL U_g1886P1975_b (.A(G1886P1975gat), .Y(G1886P1975_bgat) );
AND2XL U_g1934P2039 (.A(G1903P1793_bgat), .B(G1886P1975_bgat), .Y(G1934P2039gat) );
OR2XL U_g1949P2040 (.A(G1947P1941gat), .B(G1948P1993gat), .Y(G1949P2040gat) );
INVXL U_g1893P1972_b (.A(G1893P1972gat), .Y(G1893P1972_bgat) );
AND2XL U_g1942P2041 (.A(G1903P1793_bgat), .B(G1893P1972_bgat), .Y(G1942P2041gat) );
INVXL U_g5414P2018_b (.A(G5414P2018gat), .Y(G5414P2018_bgat) );
OR2XL U_g3964P2042 (.A(G5417P1877gat), .B(G5414P2018_bgat), .Y(G3964P2042gat) );
INVXL U_g4416P2007_b (.A(G4416P2007gat), .Y(G4416P2007_bgat) );
OR2XL U_g4425P2047 (.A(G4419P1702gat), .B(G4416P2007_bgat), .Y(G4425P2047gat) );
INVXL U_g4358P2006_b (.A(G4358P2006gat), .Y(G4358P2006_bgat) );
OR2XL U_g4367P2048 (.A(G4361P1703gat), .B(G4358P2006_bgat), .Y(G4367P2048gat) );
INVXL U_g1208P1950_b (.A(G1208P1950gat), .Y(G1208P1950_bgat) );
AND2XL U_g1256P2049 (.A(G1225P1819_bgat), .B(G1208P1950_bgat), .Y(G1256P2049gat) );
OR2XL U_g1268P2050 (.A(G1266P1954gat), .B(G1267P2003gat), .Y(G1268P2050gat) );
INVXL U_g1215P1948_b (.A(G1215P1948gat), .Y(G1215P1948_bgat) );
AND2XL U_g1261P2051 (.A(G1225P1819_bgat), .B(G1215P1948_bgat), .Y(G1261P2051gat) );
INVXL U_g4477P1825_b (.A(G4477P1825gat), .Y(G4477P1825_bgat) );
OR2XL U_g4482P2055 (.A(G4477P1825_bgat), .B(G4474P1964gat), .Y(G4482P2055gat) );
OR2XL U_g4570P2056 (.A(G1478P1731gat), .B(G4562P1965gat), .Y(G4570P2056gat) );
INVXL U_g5247P1847_b (.A(G5247P1847gat), .Y(G5247P1847_bgat) );
OR2XL U_g3536P2059 (.A(G5247P1847_bgat), .B(G5244P1966gat), .Y(G3536P2059gat) );
INVXL U_g4880P1996_b (.A(G4880P1996gat), .Y(G4880P1996_bgat) );
OR2XL U_g4889P2060 (.A(G4883P1760gat), .B(G4880P1996_bgat), .Y(G4889P2060gat) );
INVXL U_g4822P1995_b (.A(G4822P1995gat), .Y(G4822P1995_bgat) );
OR2XL U_g4831P2061 (.A(G4825P1761gat), .B(G4822P1995_bgat), .Y(G4831P2061gat) );
INVXL U_g5255P1860_b (.A(G5255P1860gat), .Y(G5255P1860_bgat) );
OR2XL U_g3541P2062 (.A(G5255P1860_bgat), .B(G5252P1976gat), .Y(G3541P2062gat) );
AND3XL U_g4074P2072 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1949P2040gat), .Y(G4074P2072gat) );
AND3XL U_g4016P2073 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1268P2050gat), .Y(G4016P2073gat) );
AND3XL U_g2347P2088 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G3850P2069gat), .Y(G2347P2088gat) );
AND3XL U_g2353P2089 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G3851P2063gat), .Y(G2353P2089gat) );
AND3XL U_g2250P2090 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G4082P2071gat), .Y(G2250P2090gat) );
AND3XL U_g2355P2091 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G3793P2065gat), .Y(G2355P2091gat) );
AND3XL U_g2349P2092 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G3792P2066gat), .Y(G2349P2092gat) );
AND3XL U_g2343P2093 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G3791P2067gat), .Y(G2343P2093gat) );
AND3XL U_g2252P2094 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G4024P2068gat), .Y(G2252P2094gat) );
AND3XL U_g1676P2095 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G3850P2069gat), .Y(G1676P2095gat) );
AND3XL U_g1682P2096 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G3851P2063gat), .Y(G1682P2096gat) );
AND3XL U_g1576P2097 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G4082P2071gat), .Y(G1576P2097gat) );
AND3XL U_g1684P2098 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G3793P2065gat), .Y(G1684P2098gat) );
AND3XL U_g1678P2099 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G3792P2066gat), .Y(G1678P2099gat) );
AND3XL U_g1672P2100 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G3791P2067gat), .Y(G1672P2100gat) );
AND3XL U_g1578P2101 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G4024P2068gat), .Y(G1578P2101gat) );
INVXL U_g5025P1987_b (.A(G5025P1987gat), .Y(G5025P1987_bgat) );
INVXL U_g5024P2036_b (.A(G5024P2036gat), .Y(G5024P2036_bgat) );
OR2XL U_g5026P2102 (.A(G5025P1987_bgat), .B(G5024P2036_bgat), .Y(G5026P2102gat) );
INVXL U_g4941P1669_b (.A(G4941P1669gat), .Y(G4941P1669_bgat) );
OR2XL U_g4946P2103 (.A(G4941P1669_bgat), .B(G4938P1989gat), .Y(G4946P2103gat) );
OR2XL U_g1944P2104 (.A(G1943P1992gat), .B(G1942P2041gat), .Y(G1944P2104gat) );
INVXL U_g5417P1877_b (.A(G5417P1877gat), .Y(G5417P1877_bgat) );
OR2XL U_g3963P2107 (.A(G5417P1877_bgat), .B(G5414P2018gat), .Y(G3963P2107gat) );
INVXL U_g5409P1998_b (.A(G5409P1998gat), .Y(G5409P1998_bgat) );
OR2XL U_g3960P2108 (.A(G5409P1998_bgat), .B(G5406P2013gat), .Y(G3960P2108gat) );
INVXL U_g4419P1702_b (.A(G4419P1702gat), .Y(G4419P1702_bgat) );
OR2XL U_g4424P2109 (.A(G4419P1702_bgat), .B(G4416P2007gat), .Y(G4424P2109gat) );
INVXL U_g4361P1703_b (.A(G4361P1703gat), .Y(G4361P1703_bgat) );
OR2XL U_g4366P2110 (.A(G4361P1703_bgat), .B(G4358P2006gat), .Y(G4366P2110gat) );
OR2XL U_g1263P2111 (.A(G1262P2002gat), .B(G1261P2051gat), .Y(G1263P2111gat) );
OR2XL U_g1258P2112 (.A(G1257P2004gat), .B(G1256P2049gat), .Y(G1258P2112gat) );
INVXL U_g4483P2010_b (.A(G4483P2010gat), .Y(G4483P2010_bgat) );
INVXL U_g4482P2055_b (.A(G4482P2055gat), .Y(G4482P2055_bgat) );
OR2XL U_g4484P2114 (.A(G4483P2010_bgat), .B(G4482P2055_bgat), .Y(G4484P2114gat) );
INVXL U_g4571P2011_b (.A(G4571P2011gat), .Y(G4571P2011_bgat) );
INVXL U_g4570P2056_b (.A(G4570P2056gat), .Y(G4570P2056_bgat) );
OR2XL U_g4572P2115 (.A(G4571P2011_bgat), .B(G4570P2056_bgat), .Y(G4572P2115gat) );
INVXL U_g5406P2013_b (.A(G5406P2013gat), .Y(G5406P2013_bgat) );
OR2XL U_g3961P2116 (.A(G5409P1998gat), .B(G5406P2013_bgat), .Y(G3961P2116gat) );
INVXL U_g4883P1760_b (.A(G4883P1760gat), .Y(G4883P1760_bgat) );
OR2XL U_g4888P2118 (.A(G4883P1760_bgat), .B(G4880P1996gat), .Y(G4888P2118gat) );
INVXL U_g4825P1761_b (.A(G4825P1761gat), .Y(G4825P1761_bgat) );
OR2XL U_g4830P2119 (.A(G4825P1761_bgat), .B(G4822P1995gat), .Y(G4830P2119gat) );
AND3XL U_g4080P2134 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1936P2105gat), .Y(G4080P2134gat) );
AND3XL U_g4077P2135 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1944P2104gat), .Y(G4077P2135gat) );
AND3XL U_g4022P2136 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1258P2112gat), .Y(G4022P2136gat) );
AND3XL U_g4019P2137 (.A(G4091P175gat), .B(G4092P176_bgat), .C(G1263P2111gat), .Y(G4019P2137gat) );
AND3XL U_g3735P2142 (.A(G3717P169gat), .B(G3724P170gat), .C(G1936P2105gat), .Y(G3735P2142gat) );
AND3XL U_g2256P2143 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G4083P2130gat), .Y(G2256P2143gat) );
AND3XL U_g2258P2144 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G4025P2129gat), .Y(G2258P2144gat) );
AND3XL U_g1582P2145 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G4083P2130gat), .Y(G1582P2145gat) );
AND3XL U_g1584P2146 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G4025P2129gat), .Y(G1584P2146gat) );
INVXL U_g5026P2102_b (.A(G5026P2102gat), .Y(G5026P2102_bgat) );
OR2XL U_g5035P2148 (.A(G5029P1668gat), .B(G5026P2102_bgat), .Y(G5035P2148gat) );
INVXL U_g4947P2038_b (.A(G4947P2038gat), .Y(G4947P2038_bgat) );
INVXL U_g4946P2103_b (.A(G4946P2103gat), .Y(G4946P2103_bgat) );
OR2XL U_g4948P2149 (.A(G4947P2038_bgat), .B(G4946P2103_bgat), .Y(G4948P2149gat) );
INVXL U_g3964P2042_b (.A(G3964P2042gat), .Y(G3964P2042_bgat) );
INVXL U_g3963P2107_b (.A(G3963P2107gat), .Y(G3963P2107_bgat) );
OR2XL U_g3965P2153 (.A(G3964P2042_bgat), .B(G3963P2107_bgat), .Y(G3965P2153gat) );
INVXL U_g3960P2108_b (.A(G3960P2108gat), .Y(G3960P2108_bgat) );
INVXL U_g3961P2116_b (.A(G3961P2116gat), .Y(G3961P2116_bgat) );
OR2XL U_g3962P2154 (.A(G3960P2108_bgat), .B(G3961P2116_bgat), .Y(G3962P2154gat) );
INVXL U_g4425P2047_b (.A(G4425P2047gat), .Y(G4425P2047_bgat) );
INVXL U_g4424P2109_b (.A(G4424P2109gat), .Y(G4424P2109_bgat) );
OR2XL U_g4426P2155 (.A(G4425P2047_bgat), .B(G4424P2109_bgat), .Y(G4426P2155gat) );
INVXL U_g4367P2048_b (.A(G4367P2048gat), .Y(G4367P2048_bgat) );
INVXL U_g4366P2110_b (.A(G4366P2110gat), .Y(G4366P2110_bgat) );
OR2XL U_g4368P2156 (.A(G4367P2048_bgat), .B(G4366P2110_bgat), .Y(G4368P2156gat) );
INVXL U_g4572P2115_b (.A(G4572P2115gat), .Y(G4572P2115_bgat) );
OR2XL U_g4581P2161 (.A(G4575P1742gat), .B(G4572P2115_bgat), .Y(G4581P2161gat) );
INVXL U_g4484P2114_b (.A(G4484P2114gat), .Y(G4484P2114_bgat) );
OR2XL U_g4493P2162 (.A(G4487P1743gat), .B(G4484P2114_bgat), .Y(G4493P2162gat) );
INVXL U_g4889P2060_b (.A(G4889P2060gat), .Y(G4889P2060_bgat) );
INVXL U_g4888P2118_b (.A(G4888P2118gat), .Y(G4888P2118_bgat) );
OR2XL U_g4890P2165 (.A(G4889P2060_bgat), .B(G4888P2118_bgat), .Y(G4890P2165gat) );
INVXL U_g4831P2061_b (.A(G4831P2061gat), .Y(G4831P2061_bgat) );
INVXL U_g4830P2119_b (.A(G4830P2119gat), .Y(G4830P2119_bgat) );
OR2XL U_g4832P2166 (.A(G4831P2061_bgat), .B(G4830P2119_bgat), .Y(G4832P2166gat) );
INVXL U_g4113P1859_b (.A(G4113P1859gat), .Y(G4113P1859_bgat) );
OR2XL U_g4096P2167 (.A(G1936P2105_bgat), .B(G4113P1859_bgat), .Y(G4096P2167gat) );
AND2XL U_g3648P2192 (.A(G4091P175_bgat), .B(G3962P2154gat), .Y(G3648P2192gat) );
AND2XL U_g3651P2193 (.A(G4091P175_bgat), .B(G3965P2153gat), .Y(G3651P2193gat) );
AND3XL U_g2262P2198 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G4084P2180gat), .Y(G2262P2198gat) );
AND3XL U_g2264P2199 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G4026P2185gat), .Y(G2264P2199gat) );
AND3XL U_g1588P2200 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G4084P2180gat), .Y(G1588P2200gat) );
AND3XL U_g1590P2201 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G4026P2185gat), .Y(G1590P2201gat) );
INVXL U_g5029P1668_b (.A(G5029P1668gat), .Y(G5029P1668_bgat) );
OR2XL U_g5034P2203 (.A(G5029P1668_bgat), .B(G5026P2102gat), .Y(G5034P2203gat) );
INVXL U_g4890P2165_b (.A(G4890P2165gat), .Y(G4890P2165_bgat) );
OR2XL U_g4899P2207 (.A(G2099P1419gat), .B(G4890P2165_bgat), .Y(G4899P2207gat) );
INVXL U_g4832P2166_b (.A(G4832P2166gat), .Y(G4832P2166_bgat) );
OR2XL U_g4841P2208 (.A(G2099P1419gat), .B(G4832P2166_bgat), .Y(G4841P2208gat) );
INVXL U_g4426P2155_b (.A(G4426P2155gat), .Y(G4426P2155_bgat) );
OR2XL U_g4435P2212 (.A(G1422P1439gat), .B(G4426P2155_bgat), .Y(G4435P2212gat) );
INVXL U_g4368P2156_b (.A(G4368P2156gat), .Y(G4368P2156_bgat) );
OR2XL U_g4377P2213 (.A(G1422P1439gat), .B(G4368P2156_bgat), .Y(G4377P2213gat) );
INVXL U_g4575P1742_b (.A(G4575P1742gat), .Y(G4575P1742_bgat) );
OR2XL U_g4580P2214 (.A(G4575P1742_bgat), .B(G4572P2115gat), .Y(G4580P2214gat) );
INVXL U_g4487P1743_b (.A(G4487P1743gat), .Y(G4487P1743_bgat) );
OR2XL U_g4492P2215 (.A(G4487P1743_bgat), .B(G4484P2114gat), .Y(G4492P2215gat) );
INVXL U_g4948P2149_b (.A(G4948P2149gat), .Y(G4948P2149_bgat) );
OR2XL U_g4957P2216 (.A(G3137P914_bgat), .B(G4948P2149_bgat), .Y(G4957P2216gat) );
AND3XL U_g2268P2251 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G4085P2232gat), .Y(G2268P2251gat) );
AND3XL U_g2274P2252 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G4086P2231gat), .Y(G2274P2252gat) );
AND3XL U_g2276P2253 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G4028P2234gat), .Y(G2276P2253gat) );
AND3XL U_g2270P2254 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G4027P2235gat), .Y(G2270P2254gat) );
AND3XL U_g1594P2255 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G4085P2232gat), .Y(G1594P2255gat) );
AND3XL U_g1600P2256 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G4086P2231gat), .Y(G1600P2256gat) );
AND3XL U_g1602P2257 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G4028P2234gat), .Y(G1602P2257gat) );
AND3XL U_g1596P2258 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G4027P2235gat), .Y(G1596P2258gat) );
INVXL U_g5035P2148_b (.A(G5035P2148gat), .Y(G5035P2148_bgat) );
INVXL U_g5034P2203_b (.A(G5034P2203gat), .Y(G5034P2203_bgat) );
OR2XL U_g5036P2259 (.A(G5035P2148_bgat), .B(G5034P2203_bgat), .Y(G5036P2259gat) );
INVXL U_g2099P1419_b (.A(G2099P1419gat), .Y(G2099P1419_bgat) );
OR2XL U_g4898P2261 (.A(G2099P1419_bgat), .B(G4890P2165gat), .Y(G4898P2261gat) );
OR2XL U_g4840P2262 (.A(G2099P1419_bgat), .B(G4832P2166gat), .Y(G4840P2262gat) );
INVXL U_g1422P1439_b (.A(G1422P1439gat), .Y(G1422P1439_bgat) );
OR2XL U_g4434P2263 (.A(G1422P1439_bgat), .B(G4426P2155gat), .Y(G4434P2263gat) );
OR2XL U_g4376P2264 (.A(G1422P1439_bgat), .B(G4368P2156gat), .Y(G4376P2264gat) );
INVXL U_g4581P2161_b (.A(G4581P2161gat), .Y(G4581P2161_bgat) );
INVXL U_g4580P2214_b (.A(G4580P2214gat), .Y(G4580P2214_bgat) );
OR2XL U_g4582P2265 (.A(G4581P2161_bgat), .B(G4580P2214_bgat), .Y(G4582P2265gat) );
INVXL U_g4493P2162_b (.A(G4493P2162gat), .Y(G4493P2162_bgat) );
INVXL U_g4492P2215_b (.A(G4492P2215gat), .Y(G4492P2215_bgat) );
OR2XL U_g4494P2266 (.A(G4493P2162_bgat), .B(G4492P2215_bgat), .Y(G4494P2266gat) );
OR2XL U_g4956P2267 (.A(G3137P914gat), .B(G4948P2149gat), .Y(G4956P2267gat) );
INVXL U_g4899P2207_b (.A(G4899P2207gat), .Y(G4899P2207_bgat) );
INVXL U_g4898P2261_b (.A(G4898P2261gat), .Y(G4898P2261_bgat) );
OR2XL U_g4900P2281 (.A(G4899P2207_bgat), .B(G4898P2261_bgat), .Y(G4900P2281gat) );
INVXL U_g4841P2208_b (.A(G4841P2208gat), .Y(G4841P2208_bgat) );
INVXL U_g4840P2262_b (.A(G4840P2262gat), .Y(G4840P2262_bgat) );
OR2XL U_g4842P2282 (.A(G4841P2208_bgat), .B(G4840P2262_bgat), .Y(G4842P2282gat) );
INVXL U_g4435P2212_b (.A(G4435P2212gat), .Y(G4435P2212_bgat) );
INVXL U_g4434P2263_b (.A(G4434P2263gat), .Y(G4434P2263_bgat) );
OR2XL U_g4436P2283 (.A(G4435P2212_bgat), .B(G4434P2263_bgat), .Y(G4436P2283gat) );
INVXL U_g4377P2213_b (.A(G4377P2213gat), .Y(G4377P2213_bgat) );
INVXL U_g4376P2264_b (.A(G4376P2264gat), .Y(G4376P2264_bgat) );
OR2XL U_g4378P2284 (.A(G4377P2213_bgat), .B(G4376P2264_bgat), .Y(G4378P2284gat) );
INVXL U_g4582P2265_b (.A(G4582P2265gat), .Y(G4582P2265_bgat) );
OR2XL U_g4591P2287 (.A(G1430P1451gat), .B(G4582P2265_bgat), .Y(G4591P2287gat) );
INVXL U_g4494P2266_b (.A(G4494P2266gat), .Y(G4494P2266_bgat) );
OR2XL U_g4503P2288 (.A(G1430P1451gat), .B(G4494P2266_bgat), .Y(G4503P2288gat) );
INVXL U_g5036P2259_b (.A(G5036P2259gat), .Y(G5036P2259_bgat) );
OR2XL U_g5045P2289 (.A(G3137P914_bgat), .B(G5036P2259_bgat), .Y(G5045P2289gat) );
INVXL U_g4957P2216_b (.A(G4957P2216gat), .Y(G4957P2216_bgat) );
INVXL U_g4956P2267_b (.A(G4956P2267gat), .Y(G4956P2267_bgat) );
OR2XL U_g4958P2290 (.A(G4957P2216_bgat), .B(G4956P2267_bgat), .Y(G4958P2290gat) );
INVXL U_g4958P2290_b (.A(G4958P2290gat), .Y(G4958P2290_bgat) );
OR2XL U_g4967P2301 (.A(G2067P1403gat), .B(G4958P2290_bgat), .Y(G4967P2301gat) );
INVXL U_g4842P2282_b (.A(G4842P2282gat), .Y(G4842P2282_bgat) );
OR2XL U_g4851P2304 (.A(G1984P1423gat), .B(G4842P2282_bgat), .Y(G4851P2304gat) );
INVXL U_g4900P2281_b (.A(G4900P2281gat), .Y(G4900P2281_bgat) );
OR2XL U_g4909P2305 (.A(G1984P1423gat), .B(G4900P2281_bgat), .Y(G4909P2305gat) );
INVXL U_g4378P2284_b (.A(G4378P2284gat), .Y(G4378P2284_bgat) );
OR2XL U_g4387P2306 (.A(G1307P1427gat), .B(G4378P2284_bgat), .Y(G4387P2306gat) );
INVXL U_g4436P2283_b (.A(G4436P2283gat), .Y(G4436P2283_bgat) );
OR2XL U_g4445P2307 (.A(G1307P1427gat), .B(G4436P2283_bgat), .Y(G4445P2307gat) );
INVXL U_g1430P1451_b (.A(G1430P1451gat), .Y(G1430P1451_bgat) );
OR2XL U_g4590P2310 (.A(G1430P1451_bgat), .B(G4582P2265gat), .Y(G4590P2310gat) );
OR2XL U_g4502P2311 (.A(G1430P1451_bgat), .B(G4494P2266gat), .Y(G4502P2311gat) );
OR2XL U_g5044P2312 (.A(G3137P914gat), .B(G5036P2259gat), .Y(G5044P2312gat) );
INVXL U_g2067P1403_b (.A(G2067P1403gat), .Y(G2067P1403_bgat) );
OR2XL U_g4966P2318 (.A(G2067P1403_bgat), .B(G4958P2290gat), .Y(G4966P2318gat) );
INVXL U_g1984P1423_b (.A(G1984P1423gat), .Y(G1984P1423_bgat) );
OR2XL U_g4850P2319 (.A(G1984P1423_bgat), .B(G4842P2282gat), .Y(G4850P2319gat) );
OR2XL U_g4908P2320 (.A(G1984P1423_bgat), .B(G4900P2281gat), .Y(G4908P2320gat) );
INVXL U_g1307P1427_b (.A(G1307P1427gat), .Y(G1307P1427_bgat) );
OR2XL U_g4386P2321 (.A(G1307P1427_bgat), .B(G4378P2284gat), .Y(G4386P2321gat) );
OR2XL U_g4444P2322 (.A(G1307P1427_bgat), .B(G4436P2283gat), .Y(G4444P2322gat) );
INVXL U_g4591P2287_b (.A(G4591P2287gat), .Y(G4591P2287_bgat) );
INVXL U_g4590P2310_b (.A(G4590P2310gat), .Y(G4590P2310_bgat) );
OR2XL U_g4592P2323 (.A(G4591P2287_bgat), .B(G4590P2310_bgat), .Y(G4592P2323gat) );
INVXL U_g4503P2288_b (.A(G4503P2288gat), .Y(G4503P2288_bgat) );
INVXL U_g4502P2311_b (.A(G4502P2311gat), .Y(G4502P2311_bgat) );
OR2XL U_g4504P2324 (.A(G4503P2288_bgat), .B(G4502P2311_bgat), .Y(G4504P2324gat) );
INVXL U_g5045P2289_b (.A(G5045P2289gat), .Y(G5045P2289_bgat) );
INVXL U_g5044P2312_b (.A(G5044P2312gat), .Y(G5044P2312_bgat) );
OR2XL U_g5046P2325 (.A(G5045P2289_bgat), .B(G5044P2312_bgat), .Y(G5046P2325gat) );
INVXL U_g4967P2301_b (.A(G4967P2301gat), .Y(G4967P2301_bgat) );
INVXL U_g4966P2318_b (.A(G4966P2318gat), .Y(G4966P2318_bgat) );
OR2XL U_g4968P2326 (.A(G4967P2301_bgat), .B(G4966P2318_bgat), .Y(G4968P2326gat) );
INVXL U_g5046P2325_b (.A(G5046P2325gat), .Y(G5046P2325_bgat) );
OR2XL U_g5055P2327 (.A(G2067P1403gat), .B(G5046P2325_bgat), .Y(G5055P2327gat) );
INVXL U_g4851P2304_b (.A(G4851P2304gat), .Y(G4851P2304_bgat) );
INVXL U_g4850P2319_b (.A(G4850P2319gat), .Y(G4850P2319_bgat) );
OR2XL U_g4852P2328 (.A(G4851P2304_bgat), .B(G4850P2319_bgat), .Y(G4852P2328gat) );
INVXL U_g4909P2305_b (.A(G4909P2305gat), .Y(G4909P2305_bgat) );
INVXL U_g4908P2320_b (.A(G4908P2320gat), .Y(G4908P2320_bgat) );
OR2XL U_g4910P2329 (.A(G4909P2305_bgat), .B(G4908P2320_bgat), .Y(G4910P2329gat) );
INVXL U_g4387P2306_b (.A(G4387P2306gat), .Y(G4387P2306_bgat) );
INVXL U_g4386P2321_b (.A(G4386P2321gat), .Y(G4386P2321_bgat) );
OR2XL U_g4388P2330 (.A(G4387P2306_bgat), .B(G4386P2321_bgat), .Y(G4388P2330gat) );
INVXL U_g4445P2307_b (.A(G4445P2307gat), .Y(G4445P2307_bgat) );
INVXL U_g4444P2322_b (.A(G4444P2322gat), .Y(G4444P2322_bgat) );
OR2XL U_g4446P2331 (.A(G4445P2307_bgat), .B(G4444P2322_bgat), .Y(G4446P2331gat) );
INVXL U_g4504P2324_b (.A(G4504P2324gat), .Y(G4504P2324_bgat) );
OR2XL U_g4513P2332 (.A(G1390P1443gat), .B(G4504P2324_bgat), .Y(G4513P2332gat) );
INVXL U_g4592P2323_b (.A(G4592P2323gat), .Y(G4592P2323_bgat) );
OR2XL U_g4601P2333 (.A(G1390P1443gat), .B(G4592P2323_bgat), .Y(G4601P2333gat) );
OR2XL U_g5054P2338 (.A(G2067P1403_bgat), .B(G5046P2325gat), .Y(G5054P2338gat) );
INVXL U_g4968P2326_b (.A(G4968P2326gat), .Y(G4968P2326_bgat) );
OR2XL U_g4977P2339 (.A(G2009P1416gat), .B(G4968P2326_bgat), .Y(G4977P2339gat) );
INVXL U_g4446P2331_b (.A(G4446P2331gat), .Y(G4446P2331_bgat) );
OR2XL U_g4455P2344 (.A(G1278P1433gat), .B(G4446P2331_bgat), .Y(G4455P2344gat) );
INVXL U_g4388P2330_b (.A(G4388P2330gat), .Y(G4388P2330_bgat) );
OR2XL U_g4397P2345 (.A(G1278P1433gat), .B(G4388P2330_bgat), .Y(G4397P2345gat) );
INVXL U_g1390P1443_b (.A(G1390P1443gat), .Y(G1390P1443_bgat) );
OR2XL U_g4512P2346 (.A(G1390P1443_bgat), .B(G4504P2324gat), .Y(G4512P2346gat) );
OR2XL U_g4600P2347 (.A(G1390P1443_bgat), .B(G4592P2323gat), .Y(G4600P2347gat) );
INVXL U_g4910P2329_b (.A(G4910P2329gat), .Y(G4910P2329_bgat) );
OR2XL U_g4919P2348 (.A(G3167P931_bgat), .B(G4910P2329_bgat), .Y(G4919P2348gat) );
INVXL U_g4852P2328_b (.A(G4852P2328gat), .Y(G4852P2328_bgat) );
OR2XL U_g4861P2349 (.A(G3167P931_bgat), .B(G4852P2328_bgat), .Y(G4861P2349gat) );
INVXL U_g5055P2327_b (.A(G5055P2327gat), .Y(G5055P2327_bgat) );
INVXL U_g5054P2338_b (.A(G5054P2338gat), .Y(G5054P2338_bgat) );
OR2XL U_g5056P2350 (.A(G5055P2327_bgat), .B(G5054P2338_bgat), .Y(G5056P2350gat) );
INVXL U_g2009P1416_b (.A(G2009P1416gat), .Y(G2009P1416_bgat) );
OR2XL U_g4976P2351 (.A(G2009P1416_bgat), .B(G4968P2326gat), .Y(G4976P2351gat) );
INVXL U_g1278P1433_b (.A(G1278P1433gat), .Y(G1278P1433_bgat) );
OR2XL U_g4454P2352 (.A(G1278P1433_bgat), .B(G4446P2331gat), .Y(G4454P2352gat) );
OR2XL U_g4396P2353 (.A(G1278P1433_bgat), .B(G4388P2330gat), .Y(G4396P2353gat) );
INVXL U_g4513P2332_b (.A(G4513P2332gat), .Y(G4513P2332_bgat) );
INVXL U_g4512P2346_b (.A(G4512P2346gat), .Y(G4512P2346_bgat) );
OR2XL U_g4514P2354 (.A(G4513P2332_bgat), .B(G4512P2346_bgat), .Y(G4514P2354gat) );
INVXL U_g4601P2333_b (.A(G4601P2333gat), .Y(G4601P2333_bgat) );
INVXL U_g4600P2347_b (.A(G4600P2347gat), .Y(G4600P2347_bgat) );
OR2XL U_g4602P2355 (.A(G4601P2333_bgat), .B(G4600P2347_bgat), .Y(G4602P2355gat) );
OR2XL U_g4918P2356 (.A(G3167P931gat), .B(G4910P2329gat), .Y(G4918P2356gat) );
OR2XL U_g4860P2357 (.A(G3167P931gat), .B(G4852P2328gat), .Y(G4860P2357gat) );
INVXL U_g5056P2350_b (.A(G5056P2350gat), .Y(G5056P2350_bgat) );
OR2XL U_g5065P2359 (.A(G2009P1416gat), .B(G5056P2350_bgat), .Y(G5065P2359gat) );
INVXL U_g4977P2339_b (.A(G4977P2339gat), .Y(G4977P2339_bgat) );
INVXL U_g4976P2351_b (.A(G4976P2351gat), .Y(G4976P2351_bgat) );
OR2XL U_g4978P2360 (.A(G4977P2339_bgat), .B(G4976P2351_bgat), .Y(G4978P2360gat) );
INVXL U_g4455P2344_b (.A(G4455P2344gat), .Y(G4455P2344_bgat) );
INVXL U_g4454P2352_b (.A(G4454P2352gat), .Y(G4454P2352_bgat) );
OR2XL U_g4456P2361 (.A(G4455P2344_bgat), .B(G4454P2352_bgat), .Y(G4456P2361gat) );
INVXL U_g4397P2345_b (.A(G4397P2345gat), .Y(G4397P2345_bgat) );
INVXL U_g4396P2353_b (.A(G4396P2353gat), .Y(G4396P2353_bgat) );
OR2XL U_g4398P2362 (.A(G4397P2345_bgat), .B(G4396P2353_bgat), .Y(G4398P2362gat) );
INVXL U_g4602P2355_b (.A(G4602P2355gat), .Y(G4602P2355_bgat) );
OR2XL U_g4611P2363 (.A(G1332P1435gat), .B(G4602P2355_bgat), .Y(G4611P2363gat) );
INVXL U_g4514P2354_b (.A(G4514P2354gat), .Y(G4514P2354_bgat) );
OR2XL U_g4523P2364 (.A(G1332P1435gat), .B(G4514P2354_bgat), .Y(G4523P2364gat) );
INVXL U_g4919P2348_b (.A(G4919P2348gat), .Y(G4919P2348_bgat) );
INVXL U_g4918P2356_b (.A(G4918P2356gat), .Y(G4918P2356_bgat) );
OR2XL U_g4920P2367 (.A(G4919P2348_bgat), .B(G4918P2356_bgat), .Y(G4920P2367gat) );
INVXL U_g4861P2349_b (.A(G4861P2349gat), .Y(G4861P2349_bgat) );
INVXL U_g4860P2357_b (.A(G4860P2357gat), .Y(G4860P2357_bgat) );
OR2XL U_g4862P2368 (.A(G4861P2349_bgat), .B(G4860P2357_bgat), .Y(G4862P2368gat) );
INVXL U_g4978P2360_b (.A(G4978P2360gat), .Y(G4978P2360_bgat) );
OR2XL U_g4987P2369 (.A(G2042P1408gat), .B(G4978P2360_bgat), .Y(G4987P2369gat) );
OR2XL U_g5064P2370 (.A(G2009P1416_bgat), .B(G5056P2350gat), .Y(G5064P2370gat) );
INVXL U_g4398P2362_b (.A(G4398P2362gat), .Y(G4398P2362_bgat) );
OR2XL U_g1488P2372 (.A(G1289P1428gat), .B(G4398P2362_bgat), .Y(G1488P2372gat) );
INVXL U_g4456P2361_b (.A(G4456P2361gat), .Y(G4456P2361_bgat) );
OR2XL U_g1493P2373 (.A(G1289P1428gat), .B(G4456P2361_bgat), .Y(G1493P2373gat) );
INVXL U_g1332P1435_b (.A(G1332P1435gat), .Y(G1332P1435_bgat) );
OR2XL U_g4610P2376 (.A(G1332P1435_bgat), .B(G4602P2355gat), .Y(G4610P2376gat) );
OR2XL U_g4522P2377 (.A(G1332P1435_bgat), .B(G4514P2354gat), .Y(G4522P2377gat) );
INVXL U_g4862P2368_b (.A(G4862P2368gat), .Y(G4862P2368_bgat) );
OR2XL U_g2165P2378 (.A(G3165P927_bgat), .B(G4862P2368_bgat), .Y(G2165P2378gat) );
INVXL U_g4920P2367_b (.A(G4920P2367gat), .Y(G4920P2367_bgat) );
OR2XL U_g2170P2379 (.A(G3165P927_bgat), .B(G4920P2367_bgat), .Y(G2170P2379gat) );
INVXL U_g2042P1408_b (.A(G2042P1408gat), .Y(G2042P1408_bgat) );
OR2XL U_g4986P2382 (.A(G2042P1408_bgat), .B(G4978P2360gat), .Y(G4986P2382gat) );
INVXL U_g5065P2359_b (.A(G5065P2359gat), .Y(G5065P2359_bgat) );
INVXL U_g5064P2370_b (.A(G5064P2370gat), .Y(G5064P2370_bgat) );
OR2XL U_g5066P2383 (.A(G5065P2359_bgat), .B(G5064P2370_bgat), .Y(G5066P2383gat) );
INVXL U_g1289P1428_b (.A(G1289P1428gat), .Y(G1289P1428_bgat) );
OR2XL U_g1487P2384 (.A(G1289P1428_bgat), .B(G4398P2362gat), .Y(G1487P2384gat) );
OR2XL U_g1492P2385 (.A(G1289P1428_bgat), .B(G4456P2361gat), .Y(G1492P2385gat) );
INVXL U_g4611P2363_b (.A(G4611P2363gat), .Y(G4611P2363_bgat) );
INVXL U_g4610P2376_b (.A(G4610P2376gat), .Y(G4610P2376_bgat) );
OR2XL U_g4612P2386 (.A(G4611P2363_bgat), .B(G4610P2376_bgat), .Y(G4612P2386gat) );
INVXL U_g4523P2364_b (.A(G4523P2364gat), .Y(G4523P2364_bgat) );
INVXL U_g4522P2377_b (.A(G4522P2377gat), .Y(G4522P2377_bgat) );
OR2XL U_g4524P2387 (.A(G4523P2364_bgat), .B(G4522P2377_bgat), .Y(G4524P2387gat) );
OR2XL U_g2164P2388 (.A(G3165P927gat), .B(G4862P2368gat), .Y(G2164P2388gat) );
OR2XL U_g2169P2389 (.A(G3165P927gat), .B(G4920P2367gat), .Y(G2169P2389gat) );
INVXL U_g5066P2383_b (.A(G5066P2383gat), .Y(G5066P2383_bgat) );
OR2XL U_g4997P2390 (.A(G2042P1408gat), .B(G5066P2383_bgat), .Y(G4997P2390gat) );
INVXL U_g4987P2369_b (.A(G4987P2369gat), .Y(G4987P2369_bgat) );
INVXL U_g4986P2382_b (.A(G4986P2382gat), .Y(G4986P2382_bgat) );
OR2XL U_g4988P2391 (.A(G4987P2369_bgat), .B(G4986P2382_bgat), .Y(G4988P2391gat) );
INVXL U_g1488P2372_b (.A(G1488P2372gat), .Y(G1488P2372_bgat) );
INVXL U_g1487P2384_b (.A(G1487P2384gat), .Y(G1487P2384_bgat) );
OR2XL U_g1489P2393 (.A(G1488P2372_bgat), .B(G1487P2384_bgat), .Y(G1489P2393gat) );
INVXL U_g1493P2373_b (.A(G1493P2373gat), .Y(G1493P2373_bgat) );
INVXL U_g1492P2385_b (.A(G1492P2385gat), .Y(G1492P2385_bgat) );
OR2XL U_g1494P2394 (.A(G1493P2373_bgat), .B(G1492P2385_bgat), .Y(G1494P2394gat) );
INVXL U_g4612P2386_b (.A(G4612P2386gat), .Y(G4612P2386_bgat) );
OR2XL U_g4543P2397 (.A(G1365P1445gat), .B(G4612P2386_bgat), .Y(G4543P2397gat) );
INVXL U_g4524P2387_b (.A(G4524P2387gat), .Y(G4524P2387_bgat) );
OR2XL U_g4533P2398 (.A(G1365P1445gat), .B(G4524P2387_bgat), .Y(G4533P2398gat) );
INVXL U_g2165P2378_b (.A(G2165P2378gat), .Y(G2165P2378_bgat) );
INVXL U_g2164P2388_b (.A(G2164P2388gat), .Y(G2164P2388_bgat) );
OR2XL U_g2166P2399 (.A(G2165P2378_bgat), .B(G2164P2388_bgat), .Y(G2166P2399gat) );
INVXL U_g2170P2379_b (.A(G2170P2379gat), .Y(G2170P2379_bgat) );
INVXL U_g2169P2389_b (.A(G2169P2389gat), .Y(G2169P2389_bgat) );
OR2XL U_g2171P2400 (.A(G2170P2379_bgat), .B(G2169P2389_bgat), .Y(G2171P2400gat) );
INVXL U_g2174P161_b (.A(G2174P161gat), .Y(G2174P161_bgat) );
AND3XL U_g2190P2401 (.A(G2174P161_bgat), .B(G2135P1673_bgat), .C(G2171P2400gat), .Y(G2190P2401gat) );
AND3XL U_g2191P2402 (.A(G2174P161_bgat), .B(G2135P1673gat), .C(G2166P2399gat), .Y(G2191P2402gat) );
INVXL U_g2160P1916_b (.A(G2160P1916gat), .Y(G2160P1916_bgat) );
AND3XL U_g2193P2403 (.A(G2174P161gat), .B(G2160P1916_bgat), .C(G2166P2399gat), .Y(G2193P2403gat) );
AND3XL U_g2192P2404 (.A(G2174P161gat), .B(G2160P1916gat), .C(G2171P2400gat), .Y(G2192P2404gat) );
INVXL U_g1497P156_b (.A(G1497P156gat), .Y(G1497P156_bgat) );
AND3XL U_g1513P2405 (.A(G1497P156_bgat), .B(G1458P1719_bgat), .C(G1494P2394gat), .Y(G1513P2405gat) );
AND3XL U_g1514P2406 (.A(G1497P156_bgat), .B(G1458P1719gat), .C(G1489P2393gat), .Y(G1514P2406gat) );
INVXL U_g1483P1895_b (.A(G1483P1895gat), .Y(G1483P1895_bgat) );
AND3XL U_g1516P2407 (.A(G1497P156gat), .B(G1483P1895_bgat), .C(G1489P2393gat), .Y(G1516P2407gat) );
AND3XL U_g1515P2408 (.A(G1497P156gat), .B(G1483P1895gat), .C(G1494P2394gat), .Y(G1515P2408gat) );
OR2XL U_g4996P2409 (.A(G2042P1408_bgat), .B(G5066P2383gat), .Y(G4996P2409gat) );
INVXL U_g4988P2391_b (.A(G4988P2391gat), .Y(G4988P2391_bgat) );
OR2XL U_g2184P2411 (.A(G2021P1306gat), .B(G4988P2391_bgat), .Y(G2184P2411gat) );
INVXL U_g1365P1445_b (.A(G1365P1445gat), .Y(G1365P1445_bgat) );
OR2XL U_g4542P2412 (.A(G1365P1445_bgat), .B(G4612P2386gat), .Y(G4542P2412gat) );
OR2XL U_g4532P2413 (.A(G1365P1445_bgat), .B(G4524P2387gat), .Y(G4532P2413gat) );
OR4XL U_g5074P2414 (.A(G2190P2401gat), .B(G2191P2402gat), .C(G2193P2403gat), .D(G2192P2404gat), .Y(G5074P2414gat) );
OR4XL U_g4620P2415 (.A(G1513P2405gat), .B(G1514P2406gat), .C(G1516P2407gat), .D(G1515P2408gat), .Y(G4620P2415gat) );
INVXL U_g4997P2390_b (.A(G4997P2390gat), .Y(G4997P2390_bgat) );
INVXL U_g4996P2409_b (.A(G4996P2409gat), .Y(G4996P2409_bgat) );
OR2XL U_g4998P2416 (.A(G4997P2390_bgat), .B(G4996P2409_bgat), .Y(G4998P2416gat) );
INVXL U_g2021P1306_b (.A(G2021P1306gat), .Y(G2021P1306_bgat) );
OR2XL U_g2183P2417 (.A(G2021P1306_bgat), .B(G4988P2391gat), .Y(G2183P2417gat) );
INVXL U_g4543P2397_b (.A(G4543P2397gat), .Y(G4543P2397_bgat) );
INVXL U_g4542P2412_b (.A(G4542P2412gat), .Y(G4542P2412_bgat) );
OR2XL U_g4544P2418 (.A(G4543P2397_bgat), .B(G4542P2412_bgat), .Y(G4544P2418gat) );
INVXL U_g4533P2398_b (.A(G4533P2398gat), .Y(G4533P2398_bgat) );
INVXL U_g4532P2413_b (.A(G4532P2413gat), .Y(G4532P2413_bgat) );
OR2XL U_g4534P2419 (.A(G4533P2398_bgat), .B(G4532P2413_bgat), .Y(G4534P2419gat) );
INVXL U_g4998P2416_b (.A(G4998P2416gat), .Y(G4998P2416_bgat) );
OR2XL U_g2187P2423 (.A(G2021P1306gat), .B(G4998P2416_bgat), .Y(G2187P2423gat) );
INVXL U_g2184P2411_b (.A(G2184P2411gat), .Y(G2184P2411_bgat) );
INVXL U_g2183P2417_b (.A(G2183P2417gat), .Y(G2183P2417_bgat) );
OR2XL U_g2185P2424 (.A(G2184P2411_bgat), .B(G2183P2417_bgat), .Y(G2185P2424gat) );
INVXL U_g4544P2418_b (.A(G4544P2418gat), .Y(G4544P2418_bgat) );
OR2XL U_g1510P2427 (.A(G1344P1449gat), .B(G4544P2418_bgat), .Y(G1510P2427gat) );
INVXL U_g4534P2419_b (.A(G4534P2419gat), .Y(G4534P2419_bgat) );
OR2XL U_g1507P2428 (.A(G1344P1449gat), .B(G4534P2419_bgat), .Y(G1507P2428gat) );
AND2XL U_g2195P2429 (.A(G2174P161gat), .B(G2185P2424gat), .Y(G2195P2429gat) );
OR2XL U_g2186P2430 (.A(G2021P1306_bgat), .B(G4998P2416gat), .Y(G2186P2430gat) );
INVXL U_g1344P1449_b (.A(G1344P1449gat), .Y(G1344P1449_bgat) );
OR2XL U_g1509P2431 (.A(G1344P1449_bgat), .B(G4544P2418gat), .Y(G1509P2431gat) );
OR2XL U_g1506P2432 (.A(G1344P1449_bgat), .B(G4534P2419gat), .Y(G1506P2432gat) );
INVXL U_g2187P2423_b (.A(G2187P2423gat), .Y(G2187P2423_bgat) );
INVXL U_g2186P2430_b (.A(G2186P2430gat), .Y(G2186P2430_bgat) );
OR2XL U_g2188P2433 (.A(G2187P2423_bgat), .B(G2186P2430_bgat), .Y(G2188P2433gat) );
INVXL U_g1510P2427_b (.A(G1510P2427gat), .Y(G1510P2427_bgat) );
INVXL U_g1509P2431_b (.A(G1509P2431gat), .Y(G1509P2431_bgat) );
OR2XL U_g1511P2434 (.A(G1510P2427_bgat), .B(G1509P2431_bgat), .Y(G1511P2434gat) );
INVXL U_g1507P2428_b (.A(G1507P2428gat), .Y(G1507P2428_bgat) );
INVXL U_g1506P2432_b (.A(G1506P2432gat), .Y(G1506P2432_bgat) );
OR2XL U_g1508P2435 (.A(G1507P2428_bgat), .B(G1506P2432_bgat), .Y(G1508P2435gat) );
AND2XL U_g1518P2436 (.A(G1497P156gat), .B(G1508P2435gat), .Y(G1518P2436gat) );
INVXL U_g2188P2433_b (.A(G2188P2433gat), .Y(G2188P2433_bgat) );
AND2XL U_g2194P2439 (.A(G2174P161_bgat), .B(G2188P2433_bgat), .Y(G2194P2439gat) );
INVXL U_g1511P2434_b (.A(G1511P2434gat), .Y(G1511P2434_bgat) );
AND2XL U_g1517P2440 (.A(G1497P156_bgat), .B(G1511P2434_bgat), .Y(G1517P2440gat) );
OR2XL U_g5077P2441 (.A(G2195P2429gat), .B(G2194P2439gat), .Y(G5077P2441gat) );
OR2XL U_g4623P2442 (.A(G1518P2436gat), .B(G1517P2440gat), .Y(G4623P2442gat) );
INVXL U_g5077P2441_b (.A(G5077P2441gat), .Y(G5077P2441_bgat) );
OR2XL U_g2196P2443 (.A(G5074P2414gat), .B(G5077P2441_bgat), .Y(G2196P2443gat) );
INVXL U_g4623P2442_b (.A(G4623P2442gat), .Y(G4623P2442_bgat) );
OR2XL U_g1519P2445 (.A(G4620P2415gat), .B(G4623P2442_bgat), .Y(G1519P2445gat) );
INVXL U_g5074P2414_b (.A(G5074P2414gat), .Y(G5074P2414_bgat) );
OR2XL U_g2197P2447 (.A(G5074P2414_bgat), .B(G5077P2441gat), .Y(G2197P2447gat) );
INVXL U_g4620P2415_b (.A(G4620P2415gat), .Y(G4620P2415_bgat) );
OR2XL U_g1520P2448 (.A(G4620P2415_bgat), .B(G4623P2442gat), .Y(G1520P2448gat) );
INVXL U_g2196P2443_b (.A(G2196P2443gat), .Y(G2196P2443_bgat) );
INVXL U_g2197P2447_b (.A(G2197P2447gat), .Y(G2197P2447_bgat) );
OR2XL U_g2198P2449 (.A(G2196P2443_bgat), .B(G2197P2447_bgat), .Y(G2198P2449gat) );
INVXL U_g1519P2445_b (.A(G1519P2445gat), .Y(G1519P2445_bgat) );
INVXL U_g1520P2448_b (.A(G1520P2448gat), .Y(G1520P2448_bgat) );
OR2XL U_g1521P2450 (.A(G1519P2445_bgat), .B(G1520P2448_bgat), .Y(G1521P2450gat) );
INVXL U_g2198P2449_b (.A(G2198P2449gat), .Y(G2198P2449_bgat) );
AND2XL U_g3652P2457 (.A(G4091P175gat), .B(G2198P2449_bgat), .Y(G3652P2457gat) );
INVXL U_g1521P2450_b (.A(G1521P2450gat), .Y(G1521P2450_bgat) );
AND2XL U_g3649P2458 (.A(G4091P175gat), .B(G1521P2450_bgat), .Y(G3649P2458gat) );
OR2XL U_g3657P2459 (.A(G3648P2192gat), .B(G3649P2458gat), .Y(G3657P2459gat) );
OR2XL U_g3658P2460 (.A(G3651P2193gat), .B(G3652P2457gat), .Y(G3658P2460gat) );
AND2XL U_g3636P2461 (.A(G4092P176_bgat), .B(G3657P2459gat), .Y(G3636P2461gat) );
AND2XL U_g3642P2462 (.A(G4092P176_bgat), .B(G3657P2459gat), .Y(G3642P2462gat) );
AND2XL U_g3639P2463 (.A(G4092P176_bgat), .B(G3658P2460gat), .Y(G3639P2463gat) );
AND2XL U_g3645P2464 (.A(G4092P176_bgat), .B(G3658P2460gat), .Y(G3645P2464gat) );
OR2XL U_g3655P2465 (.A(G3643P634gat), .B(G3642P2462gat), .Y(G3655P2465gat) );
OR2XL U_g3653P2466 (.A(G3637P635gat), .B(G3636P2461gat), .Y(G3653P2466gat) );
OR2XL U_g3656P2467 (.A(G3646P636gat), .B(G3645P2464gat), .Y(G3656P2467gat) );
OR2XL U_g3654P2468 (.A(G3640P637gat), .B(G3639P2463gat), .Y(G3654P2468gat) );
AND3XL U_g2328P2473 (.A(G1691P159_bgat), .B(G1694P160_bgat), .C(G3654P2468gat), .Y(G2328P2473gat) );
AND3XL U_g2330P2474 (.A(G1691P159gat), .B(G1694P160_bgat), .C(G3653P2466gat), .Y(G2330P2474gat) );
AND3XL U_g1657P2475 (.A(G1689P157_bgat), .B(G1690P158_bgat), .C(G3654P2468gat), .Y(G1657P2475gat) );
AND3XL U_g1659P2476 (.A(G1689P157gat), .B(G1690P158_bgat), .C(G3653P2466gat), .Y(G1659P2476gat) );
OR4XL U_g1662P2477 (.A(G1661P601gat), .B(G1660P799gat), .C(G1657P2475gat), .D(G1659P2476gat), .Y(G1662P2477gat) );
OR4XL U_g2333P2478 (.A(G2332P602gat), .B(G2331P798gat), .C(G2328P2473gat), .D(G2330P2474gat), .Y(G2333P2478gat) );

endmodule
