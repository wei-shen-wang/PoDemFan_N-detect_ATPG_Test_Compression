module C880 ( G1GAT_0_gat, G8GAT_1_gat, G13GAT_2_gat, G17GAT_3_gat, G26GAT_4_gat, G29GAT_5_gat, G36GAT_6_gat, G42GAT_7_gat, G51GAT_8_gat, G55GAT_9_gat, G59GAT_10_gat, G68GAT_11_gat, G72GAT_12_gat, G73GAT_13_gat, G74GAT_14_gat, G75GAT_15_gat, G80GAT_16_gat, G85GAT_17_gat, G86GAT_18_gat, G87GAT_19_gat, G88GAT_20_gat, G89GAT_21_gat, G90GAT_22_gat, G91GAT_23_gat, G96GAT_24_gat, G101GAT_25_gat, G106GAT_26_gat, G111GAT_27_gat, G116GAT_28_gat, G121GAT_29_gat, G126GAT_30_gat, G130GAT_31_gat, G135GAT_32_gat, G138GAT_33_gat, G143GAT_34_gat, G146GAT_35_gat, G149GAT_36_gat, G152GAT_37_gat, G153GAT_38_gat, G156GAT_39_gat, G159GAT_40_gat, G165GAT_41_gat, G171GAT_42_gat, G177GAT_43_gat, G183GAT_44_gat, G189GAT_45_gat, G195GAT_46_gat, G201GAT_47_gat, G207GAT_48_gat, G210GAT_49_gat, G219GAT_50_gat, G228GAT_51_gat, G237GAT_52_gat, G246GAT_53_gat, G255GAT_54_gat, G259GAT_55_gat, G260GAT_56_gat, G261GAT_57_gat, G267GAT_58_gat, G268GAT_59_gat, G388GAT_133_gat, G389GAT_132_gat, G390GAT_131_gat, G391GAT_124_gat, G418GAT_168_gat, G419GAT_164_gat, G420GAT_158_gat, G421GAT_162_gat, G422GAT_161_gat, G423GAT_155_gat, G446GAT_183_gat, G447GAT_182_gat, G448GAT_179_gat, G449GAT_176_gat, G450GAT_173_gat, G767GAT_349_gat, G768GAT_334_gat, G850GAT_404_gat, G863GAT_424_gat, G864GAT_423_gat, G865GAT_422_gat, G866GAT_426_gat, G874GAT_433_gat, G878GAT_442_gat, G879GAT_441_gat, G880GAT_440_gat);

input G1GAT_0_gat;
input G8GAT_1_gat;
input G13GAT_2_gat;
input G17GAT_3_gat;
input G26GAT_4_gat;
input G29GAT_5_gat;
input G36GAT_6_gat;
input G42GAT_7_gat;
input G51GAT_8_gat;
input G55GAT_9_gat;
input G59GAT_10_gat;
input G68GAT_11_gat;
input G72GAT_12_gat;
input G73GAT_13_gat;
input G74GAT_14_gat;
input G75GAT_15_gat;
input G80GAT_16_gat;
input G85GAT_17_gat;
input G86GAT_18_gat;
input G87GAT_19_gat;
input G88GAT_20_gat;
input G89GAT_21_gat;
input G90GAT_22_gat;
input G91GAT_23_gat;
input G96GAT_24_gat;
input G101GAT_25_gat;
input G106GAT_26_gat;
input G111GAT_27_gat;
input G116GAT_28_gat;
input G121GAT_29_gat;
input G126GAT_30_gat;
input G130GAT_31_gat;
input G135GAT_32_gat;
input G138GAT_33_gat;
input G143GAT_34_gat;
input G146GAT_35_gat;
input G149GAT_36_gat;
input G152GAT_37_gat;
input G153GAT_38_gat;
input G156GAT_39_gat;
input G159GAT_40_gat;
input G165GAT_41_gat;
input G171GAT_42_gat;
input G177GAT_43_gat;
input G183GAT_44_gat;
input G189GAT_45_gat;
input G195GAT_46_gat;
input G201GAT_47_gat;
input G207GAT_48_gat;
input G210GAT_49_gat;
input G219GAT_50_gat;
input G228GAT_51_gat;
input G237GAT_52_gat;
input G246GAT_53_gat;
input G255GAT_54_gat;
input G259GAT_55_gat;
input G260GAT_56_gat;
input G261GAT_57_gat;
input G267GAT_58_gat;
input G268GAT_59_gat;

output G388GAT_133_gat;
output G389GAT_132_gat;
output G390GAT_131_gat;
output G391GAT_124_gat;
output G418GAT_168_gat;
output G419GAT_164_gat;
output G420GAT_158_gat;
output G421GAT_162_gat;
output G422GAT_161_gat;
output G423GAT_155_gat;
output G446GAT_183_gat;
output G447GAT_182_gat;
output G448GAT_179_gat;
output G449GAT_176_gat;
output G450GAT_173_gat;
output G767GAT_349_gat;
output G768GAT_334_gat;
output G850GAT_404_gat;
output G863GAT_424_gat;
output G864GAT_423_gat;
output G865GAT_422_gat;
output G866GAT_426_gat;
output G874GAT_433_gat;
output G878GAT_442_gat;
output G879GAT_441_gat;
output G880GAT_440_gat;

BUFX20 U_g1 (.A(G268GAT_59_gat), .Y(G310GAT_60_gat) );
AND2XL U_g2 (.A(G267GAT_58_gat), .B(G255GAT_54_gat), .Y(G341GAT_61_gat) );
AND2XL U_g3 (.A(G260GAT_56_gat), .B(G255GAT_54_gat), .Y(G339GAT_62_gat) );
AND2XL U_g4 (.A(G259GAT_55_gat), .B(G255GAT_54_gat), .Y(G337GAT_63_gat) );
AND2XL U_g5 (.A(G201GAT_47_ngat), .B(G195GAT_46_ngat), .Y(G331GAT_64_gat) );
AND2XL U_g6 (.A(G201GAT_47_gat), .B(G195GAT_46_gat), .Y(G330GAT_65_gat) );
AND2XL U_g7 (.A(G189GAT_45_ngat), .B(G183GAT_44_ngat), .Y(G329GAT_66_gat) );
AND2XL U_g8 (.A(G189GAT_45_gat), .B(G183GAT_44_gat), .Y(G328GAT_67_gat) );
AND2XL U_g9 (.A(G177GAT_43_ngat), .B(G171GAT_42_ngat), .Y(G327GAT_68_gat) );
AND2XL U_g10 (.A(G177GAT_43_gat), .B(G171GAT_42_gat), .Y(G326GAT_69_gat) );
AND2XL U_g11 (.A(G165GAT_41_ngat), .B(G159GAT_40_ngat), .Y(G325GAT_70_gat) );
AND2XL U_g12 (.A(G165GAT_41_gat), .B(G159GAT_40_gat), .Y(G324GAT_71_gat) );
AND2XL U_g13 (.A(G138GAT_33_gat), .B(G152GAT_37_gat), .Y(G318GAT_72_gat) );
AND2XL U_g14 (.A(G121GAT_29_gat), .B(G210GAT_49_gat), .Y(G340GAT_73_gat) );
AND2XL U_g15 (.A(G126GAT_30_ngat), .B(G121GAT_29_ngat), .Y(G308GAT_74_gat) );
AND2XL U_g16 (.A(G126GAT_30_gat), .B(G121GAT_29_gat), .Y(G307GAT_75_gat) );
AND2XL U_g17 (.A(G116GAT_28_gat), .B(G210GAT_49_gat), .Y(G338GAT_76_gat) );
AND2XL U_g18 (.A(G111GAT_27_gat), .B(G210GAT_49_gat), .Y(G336GAT_77_gat) );
AND2XL U_g19 (.A(G116GAT_28_ngat), .B(G111GAT_27_ngat), .Y(G306GAT_78_gat) );
AND2XL U_g20 (.A(G116GAT_28_gat), .B(G111GAT_27_gat), .Y(G305GAT_79_gat) );
AND2XL U_g21 (.A(G106GAT_26_gat), .B(G210GAT_49_gat), .Y(G335GAT_80_gat) );
AND2XL U_g22 (.A(G101GAT_25_gat), .B(G210GAT_49_gat), .Y(G334GAT_81_gat) );
AND2XL U_g23 (.A(G106GAT_26_ngat), .B(G101GAT_25_ngat), .Y(G304GAT_82_gat) );
AND2XL U_g24 (.A(G106GAT_26_gat), .B(G101GAT_25_gat), .Y(G303GAT_83_gat) );
AND2XL U_g25 (.A(G96GAT_24_gat), .B(G210GAT_49_gat), .Y(G333GAT_84_gat) );
AND2XL U_g26 (.A(G91GAT_23_gat), .B(G210GAT_49_gat), .Y(G332GAT_85_gat) );
AND2XL U_g27 (.A(G96GAT_24_ngat), .B(G91GAT_23_ngat), .Y(G302GAT_86_gat) );
AND2XL U_g28 (.A(G96GAT_24_gat), .B(G91GAT_23_gat), .Y(G301GAT_87_gat) );
AND2XL U_g29 (.A(G88GAT_20_ngat), .B(G87GAT_19_ngat), .Y(G298GAT_88_gat) );
AND2XL U_g30 (.A(G86GAT_18_gat), .B(G85GAT_17_gat), .Y(G297GAT_89_gat) );
AND2XL U_g31 (.A(G156GAT_39_gat), .B(G59GAT_10_gat), .Y(G319GAT_90_gat) );
AND3XL U_g32 (.A(G80GAT_16_gat), .B(G75GAT_15_gat), .C(G59GAT_10_gat), .Y(G293GAT_91_gat) );
AND3XL U_g33 (.A(G74GAT_14_gat), .B(G68GAT_11_gat), .C(G59GAT_10_gat), .Y(G286GAT_92_gat) );
AND2XL U_g34 (.A(G138GAT_33_gat), .B(G51GAT_8_gat), .Y(G316GAT_93_gat) );
AND3XL U_g35 (.A(G42GAT_7_gat), .B(G75GAT_15_gat), .C(G59GAT_10_gat), .Y(G294GAT_94_gat) );
AND4XL U_g36 (.A(G72GAT_12_gat), .B(G68GAT_11_gat), .C(G42GAT_7_gat), .D(G59GAT_10_gat), .Y(G284GAT_95_gat) );
AND3XL U_g37 (.A(G42GAT_7_gat), .B(G36GAT_6_gat), .C(G59GAT_10_gat), .Y(G296GAT_96_gat) );
AND3XL U_g38 (.A(G80GAT_16_gat), .B(G36GAT_6_gat), .C(G59GAT_10_gat), .Y(G295GAT_97_gat) );
AND3XL U_g39 (.A(G42GAT_7_gat), .B(G36GAT_6_gat), .C(G29GAT_5_gat), .Y(G292GAT_98_gat) );
AND3XL U_g40 (.A(G80GAT_16_gat), .B(G36GAT_6_gat), .C(G29GAT_5_gat), .Y(G291GAT_99_gat) );
AND3XL U_g41 (.A(G42GAT_7_gat), .B(G75GAT_15_gat), .C(G29GAT_5_gat), .Y(G290GAT_100_gat) );
AND3XL U_g42 (.A(G80GAT_16_gat), .B(G75GAT_15_gat), .C(G29GAT_5_gat), .Y(G287GAT_101_gat) );
AND2XL U_g43 (.A(G68GAT_11_gat), .B(G29GAT_5_gat), .Y(G285GAT_102_gat) );
AND3XL U_g44 (.A(G42GAT_7_gat), .B(G36GAT_6_gat), .C(G29GAT_5_gat), .Y(G273GAT_103_gat) );
AND2XL U_g45 (.A(G42GAT_7_gat), .B(G17GAT_3_gat), .Y(G323GAT_104_gat) );
AND2XL U_g46 (.A(G42GAT_7_ngat), .B(G17GAT_3_ngat), .Y(G322GAT_105_gat) );
AND2XL U_g47 (.A(G138GAT_33_gat), .B(G17GAT_3_gat), .Y(G317GAT_106_gat) );
AND2XL U_g48 (.A(G138GAT_33_gat), .B(G8GAT_1_gat), .Y(G309GAT_107_gat) );
AND4XL U_g49 (.A(G55GAT_9_gat), .B(G13GAT_2_gat), .C(G8GAT_1_gat), .D(G1GAT_0_gat), .Y(G280GAT_108_gat) );
AND4XL U_g50 (.A(G17GAT_3_gat), .B(G51GAT_8_gat), .C(G8GAT_1_gat), .D(G1GAT_0_gat), .Y(G279GAT_109_gat) );
AND3XL U_g51 (.A(G51GAT_8_gat), .B(G26GAT_4_gat), .C(G1GAT_0_gat), .Y(G276GAT_110_gat) );
AND4XL U_g52 (.A(G17GAT_3_gat), .B(G13GAT_2_gat), .C(G26GAT_4_gat), .D(G1GAT_0_gat), .Y(G270GAT_111_gat) );
AND4XL U_g53 (.A(G17GAT_3_gat), .B(G13GAT_2_gat), .C(G8GAT_1_gat), .D(G1GAT_0_gat), .Y(G269GAT_112_gat) );
BUFX20 U_g54 (.A(G310GAT_60_gat), .Y(G369GAT_113_gat) );
AND2XL U_g55 (.A(G331GAT_64_gat), .B(G330GAT_65_gat), .Y(G385GAT_114_gat) );
AND2XL U_g56 (.A(G329GAT_66_gat), .B(G328GAT_67_gat), .Y(G382GAT_115_gat) );
AND2XL U_g57 (.A(G327GAT_68_gat), .B(G326GAT_69_gat), .Y(G379GAT_116_gat) );
AND2XL U_g58 (.A(G325GAT_70_gat), .B(G324GAT_71_gat), .Y(G376GAT_117_gat) );
AND2XL U_g59 (.A(G308GAT_74_gat), .B(G307GAT_75_gat), .Y(G366GAT_118_gat) );
AND2XL U_g60 (.A(G306GAT_78_gat), .B(G305GAT_79_gat), .Y(G363GAT_119_gat) );
AND2XL U_g61 (.A(G304GAT_82_gat), .B(G303GAT_83_gat), .Y(G360GAT_120_gat) );
AND2XL U_g62 (.A(G302GAT_86_gat), .B(G301GAT_87_gat), .Y(G357GAT_121_gat) );
AND2XL U_g63 (.A(G298GAT_88_gat), .B(G90GAT_22_gat), .Y(G356GAT_122_gat) );
AND2XL U_g64 (.A(G298GAT_88_gat), .B(G89GAT_21_gat), .Y(G355GAT_123_gat) );
BUFX20 U_g65 (.A(G297GAT_89_gat), .Y(G391GAT_124_gat) );
BUFX20 U_g66 (.A(G293GAT_91_gat), .Y(G351GAT_125_gat) );
AND2XL U_g67 (.A(G286GAT_92_ngat), .B(G280GAT_108_ngat), .Y(G350GAT_126_gat) );
BUFX20 U_g68 (.A(G294GAT_94_gat), .Y(G352GAT_127_gat) );
AND2XL U_g69 (.A(G284GAT_95_ngat), .B(G280GAT_108_ngat), .Y(G348GAT_128_gat) );
BUFX20 U_g70 (.A(G296GAT_96_gat), .Y(G354GAT_129_gat) );
BUFX20 U_g71 (.A(G295GAT_97_gat), .Y(G353GAT_130_gat) );
BUFX20 U_g72 (.A(G292GAT_98_gat), .Y(G390GAT_131_gat) );
BUFX20 U_g73 (.A(G291GAT_99_gat), .Y(G389GAT_132_gat) );
BUFX20 U_g74 (.A(G290GAT_100_gat), .Y(G388GAT_133_gat) );
AND2XL U_g75 (.A(G285GAT_102_ngat), .B(G280GAT_108_ngat), .Y(G349GAT_134_gat) );
BUFX20 U_g76 (.A(G273GAT_103_gat), .Y(G343GAT_135_gat) );
AND2XL U_g77 (.A(G273GAT_103_ngat), .B(G270GAT_111_ngat), .Y(G344GAT_136_gat) );
AND2XL U_g78 (.A(G323GAT_104_ngat), .B(G322GAT_105_ngat), .Y(G375GAT_137_gat) );
BUFX20 U_g79 (.A(G279GAT_109_gat), .Y(G347GAT_138_gat) );
BUFX20 U_g80 (.A(G276GAT_110_gat), .Y(G345GAT_139_gat) );
BUFX20 U_g81 (.A(G276GAT_110_gat), .Y(G346GAT_140_gat) );
BUFX20 U_g82 (.A(G269GAT_112_gat), .Y(G342GAT_141_gat) );
AND2XL U_g83 (.A(G369GAT_113_gat), .B(G210GAT_49_gat), .Y(G417GAT_142_gat) );
BUFX20 U_g84 (.A(G385GAT_114_gat), .Y(G415GAT_143_gat) );
AND2XL U_g85 (.A(G385GAT_114_gat), .B(G382GAT_115_gat), .Y(G416GAT_144_gat) );
BUFX20 U_g86 (.A(G382GAT_115_gat), .Y(G414GAT_145_gat) );
BUFX20 U_g87 (.A(G379GAT_116_gat), .Y(G412GAT_146_gat) );
AND2XL U_g88 (.A(G379GAT_116_gat), .B(G376GAT_117_gat), .Y(G413GAT_147_gat) );
BUFX20 U_g89 (.A(G376GAT_117_gat), .Y(G411GAT_148_gat) );
BUFX20 U_g90 (.A(G366GAT_118_gat), .Y(G408GAT_149_gat) );
AND2XL U_g91 (.A(G366GAT_118_gat), .B(G363GAT_119_gat), .Y(G409GAT_150_gat) );
BUFX20 U_g92 (.A(G363GAT_119_gat), .Y(G407GAT_151_gat) );
BUFX20 U_g93 (.A(G360GAT_120_gat), .Y(G405GAT_152_gat) );
AND2XL U_g94 (.A(G360GAT_120_gat), .B(G357GAT_121_gat), .Y(G406GAT_153_gat) );
BUFX20 U_g95 (.A(G357GAT_121_gat), .Y(G404GAT_154_gat) );
BUFX20 U_g96 (.A(G356GAT_122_gat), .Y(G423GAT_155_gat) );
BUFX20 U_g97 (.A(G355GAT_123_gat), .Y(G403GAT_156_gat) );
AND2XL U_g98 (.A(G73GAT_13_gat), .B(G348GAT_128_gat), .Y(G400GAT_157_gat) );
BUFX20 U_g99 (.A(G351GAT_125_gat), .Y(G420GAT_158_gat) );
BUFX20 U_g100 (.A(G350GAT_126_gat), .Y(G402GAT_159_gat) );
AND2XL U_g101 (.A(G352GAT_127_gat), .B(G347GAT_138_gat), .Y(G410GAT_160_gat) );
BUFX20 U_g102 (.A(G354GAT_129_gat), .Y(G422GAT_161_gat) );
BUFX20 U_g103 (.A(G353GAT_130_gat), .Y(G421GAT_162_gat) );
BUFX20 U_g104 (.A(G349GAT_134_gat), .Y(G401GAT_163_gat) );
BUFX20 U_g105 (.A(G344GAT_136_gat), .Y(G419GAT_164_gat) );
BUFX20 U_g106 (.A(G345GAT_139_gat), .Y(G393GAT_165_gat) );
BUFX20 U_g107 (.A(G346GAT_140_gat), .Y(G399GAT_166_gat) );
AND2XL U_g108 (.A(G343GAT_135_ngat), .B(G270GAT_111_ngat), .Y(G392GAT_167_gat) );
BUFX20 U_g109 (.A(G342GAT_141_gat), .Y(G418GAT_168_gat) );
AND2XL U_g110 (.A(G415GAT_143_gat), .B(G414GAT_145_gat), .Y(G445GAT_169_gat) );
AND2XL U_g111 (.A(G412GAT_146_gat), .B(G411GAT_148_gat), .Y(G444GAT_170_gat) );
AND2XL U_g112 (.A(G408GAT_149_gat), .B(G407GAT_151_gat), .Y(G426GAT_171_gat) );
AND2XL U_g113 (.A(G405GAT_152_gat), .B(G404GAT_154_gat), .Y(G425GAT_172_gat) );
BUFX20 U_g114 (.A(G403GAT_156_gat), .Y(G450GAT_173_gat) );
BUFX20 U_g115 (.A(G400GAT_157_gat), .Y(G424GAT_174_gat) );
AND4XL U_g116 (.A(G393GAT_165_gat), .B(G156GAT_39_gat), .C(G59GAT_10_gat), .D(G375GAT_137_gat), .Y(G442GAT_175_gat) );
BUFX20 U_g117 (.A(G402GAT_159_gat), .Y(G449GAT_176_gat) );
AND3XL U_g118 (.A(G55GAT_9_gat), .B(G287GAT_101_gat), .C(G393GAT_165_gat), .Y(G437GAT_177_gat) );
AND3XL U_g119 (.A(G55GAT_9_gat), .B(G393GAT_165_gat), .C(G319GAT_90_gat), .Y(G427GAT_178_gat) );
BUFX20 U_g120 (.A(G401GAT_163_gat), .Y(G448GAT_179_gat) );
AND3XL U_g121 (.A(G17GAT_3_gat), .B(G319GAT_90_gat), .C(G393GAT_165_gat), .Y(G443GAT_180_gat) );
AND3XL U_g122 (.A(G287GAT_101_gat), .B(G17GAT_3_gat), .C(G393GAT_165_gat), .Y(G432GAT_181_gat) );
BUFX20 U_g123 (.A(G399GAT_166_gat), .Y(G447GAT_182_gat) );
BUFX20 U_g124 (.A(G392GAT_167_gat), .Y(G446GAT_183_gat) );
AND2XL U_g125 (.A(G437GAT_177_ngat), .B(G369GAT_113_ngat), .Y(G488GAT_184_gat) );
AND2XL U_g126 (.A(G437GAT_177_ngat), .B(G369GAT_113_ngat), .Y(G489GAT_185_gat) );
AND2XL U_g127 (.A(G437GAT_177_ngat), .B(G369GAT_113_ngat), .Y(G490GAT_186_gat) );
AND2XL U_g128 (.A(G437GAT_177_ngat), .B(G369GAT_113_ngat), .Y(G491GAT_187_gat) );
AND2XL U_g129 (.A(G432GAT_181_gat), .B(G310GAT_60_gat), .Y(G476GAT_188_gat) );
AND2XL U_g130 (.A(G432GAT_181_gat), .B(G310GAT_60_gat), .Y(G478GAT_189_gat) );
AND2XL U_g131 (.A(G432GAT_181_gat), .B(G310GAT_60_gat), .Y(G480GAT_190_gat) );
AND2XL U_g132 (.A(G432GAT_181_gat), .B(G310GAT_60_gat), .Y(G482GAT_191_gat) );
AND2XL U_g133 (.A(G445GAT_169_ngat), .B(G416GAT_144_ngat), .Y(G495GAT_192_gat) );
AND2XL U_g134 (.A(G444GAT_170_ngat), .B(G413GAT_147_ngat), .Y(G492GAT_193_gat) );
AND2XL U_g135 (.A(G427GAT_178_gat), .B(G153GAT_38_gat), .Y(G481GAT_194_gat) );
AND2XL U_g136 (.A(G427GAT_178_gat), .B(G149GAT_36_gat), .Y(G479GAT_195_gat) );
AND2XL U_g137 (.A(G427GAT_178_gat), .B(G146GAT_35_gat), .Y(G477GAT_196_gat) );
AND2XL U_g138 (.A(G427GAT_178_gat), .B(G143GAT_34_gat), .Y(G475GAT_197_gat) );
AND2XL U_g139 (.A(G426GAT_171_ngat), .B(G409GAT_150_ngat), .Y(G463GAT_198_gat) );
AND2XL U_g140 (.A(G425GAT_172_ngat), .B(G406GAT_153_ngat), .Y(G460GAT_199_gat) );
BUFX20 U_g141 (.A(G424GAT_174_gat), .Y(G451GAT_200_gat) );
AND2XL U_g142 (.A(G410GAT_160_gat), .B(G442GAT_175_gat), .Y(G466GAT_201_gat) );
AND2XL U_g143 (.A(G1GAT_0_gat), .B(G443GAT_180_gat), .Y(G483GAT_202_gat) );
AND2XL U_g144 (.A(G476GAT_188_ngat), .B(G475GAT_197_ngat), .Y(G503GAT_203_gat) );
AND2XL U_g145 (.A(G478GAT_189_ngat), .B(G477GAT_196_ngat), .Y(G505GAT_204_gat) );
AND2XL U_g146 (.A(G480GAT_190_ngat), .B(G479GAT_195_ngat), .Y(G507GAT_205_gat) );
AND2XL U_g147 (.A(G482GAT_191_ngat), .B(G481GAT_194_ngat), .Y(G509GAT_206_gat) );
AND2XL U_g148 (.A(G207GAT_48_ngat), .B(G495GAT_192_ngat), .Y(G521GAT_207_gat) );
AND2XL U_g149 (.A(G207GAT_48_gat), .B(G495GAT_192_gat), .Y(G520GAT_208_gat) );
AND2XL U_g150 (.A(G201GAT_47_gat), .B(G451GAT_200_gat), .Y(G529GAT_209_gat) );
AND2XL U_g151 (.A(G195GAT_46_gat), .B(G451GAT_200_gat), .Y(G528GAT_210_gat) );
AND2XL U_g152 (.A(G189GAT_45_gat), .B(G451GAT_200_gat), .Y(G527GAT_211_gat) );
AND2XL U_g153 (.A(G183GAT_44_gat), .B(G451GAT_200_gat), .Y(G526GAT_212_gat) );
AND2XL U_g154 (.A(G177GAT_43_gat), .B(G451GAT_200_gat), .Y(G525GAT_213_gat) );
AND2XL U_g155 (.A(G171GAT_42_gat), .B(G451GAT_200_gat), .Y(G524GAT_214_gat) );
AND2XL U_g156 (.A(G165GAT_41_gat), .B(G451GAT_200_gat), .Y(G523GAT_215_gat) );
AND2XL U_g157 (.A(G159GAT_40_gat), .B(G451GAT_200_gat), .Y(G522GAT_216_gat) );
AND2XL U_g158 (.A(G483GAT_202_gat), .B(G153GAT_38_gat), .Y(G516GAT_217_gat) );
AND2XL U_g159 (.A(G483GAT_202_gat), .B(G149GAT_36_gat), .Y(G514GAT_218_gat) );
AND2XL U_g160 (.A(G483GAT_202_gat), .B(G146GAT_35_gat), .Y(G512GAT_219_gat) );
AND2XL U_g161 (.A(G483GAT_202_gat), .B(G143GAT_34_gat), .Y(G510GAT_220_gat) );
AND2XL U_g162 (.A(G135GAT_32_ngat), .B(G463GAT_198_ngat), .Y(G501GAT_221_gat) );
AND2XL U_g163 (.A(G135GAT_32_gat), .B(G463GAT_198_gat), .Y(G500GAT_222_gat) );
AND2XL U_g164 (.A(G492GAT_193_ngat), .B(G130GAT_31_ngat), .Y(G519GAT_223_gat) );
AND2XL U_g165 (.A(G492GAT_193_gat), .B(G130GAT_31_gat), .Y(G518GAT_224_gat) );
AND2XL U_g166 (.A(G460GAT_199_ngat), .B(G130GAT_31_ngat), .Y(G499GAT_225_gat) );
AND2XL U_g167 (.A(G460GAT_199_gat), .B(G130GAT_31_gat), .Y(G498GAT_226_gat) );
AND2XL U_g168 (.A(G466GAT_201_gat), .B(G126GAT_30_gat), .Y(G517GAT_227_gat) );
AND2XL U_g169 (.A(G466GAT_201_gat), .B(G121GAT_29_gat), .Y(G515GAT_228_gat) );
AND2XL U_g170 (.A(G466GAT_201_gat), .B(G116GAT_28_gat), .Y(G513GAT_229_gat) );
AND2XL U_g171 (.A(G466GAT_201_gat), .B(G111GAT_27_gat), .Y(G511GAT_230_gat) );
AND2XL U_g172 (.A(G466GAT_201_gat), .B(G106GAT_26_gat), .Y(G508GAT_231_gat) );
AND2XL U_g173 (.A(G466GAT_201_gat), .B(G101GAT_25_gat), .Y(G506GAT_232_gat) );
AND2XL U_g174 (.A(G466GAT_201_gat), .B(G96GAT_24_gat), .Y(G504GAT_233_gat) );
AND2XL U_g175 (.A(G466GAT_201_gat), .B(G91GAT_23_gat), .Y(G502GAT_234_gat) );
AND2XL U_g176 (.A(G521GAT_207_gat), .B(G520GAT_208_gat), .Y(G547GAT_235_gat) );
AND2XL U_g177 (.A(G517GAT_227_ngat), .B(G516GAT_217_ngat), .Y(G543GAT_236_gat) );
AND2XL U_g178 (.A(G515GAT_228_ngat), .B(G514GAT_218_ngat), .Y(G542GAT_237_gat) );
AND2XL U_g179 (.A(G513GAT_229_ngat), .B(G512GAT_219_ngat), .Y(G541GAT_238_gat) );
AND2XL U_g180 (.A(G511GAT_230_ngat), .B(G510GAT_220_ngat), .Y(G540GAT_239_gat) );
AND2XL U_g181 (.A(G508GAT_231_ngat), .B(G318GAT_72_ngat), .Y(G539GAT_240_gat) );
AND2XL U_g182 (.A(G501GAT_221_gat), .B(G500GAT_222_gat), .Y(G533GAT_241_gat) );
AND2XL U_g183 (.A(G519GAT_223_gat), .B(G518GAT_224_gat), .Y(G544GAT_242_gat) );
AND2XL U_g184 (.A(G499GAT_225_gat), .B(G498GAT_226_gat), .Y(G530GAT_243_gat) );
AND2XL U_g185 (.A(G504GAT_233_ngat), .B(G316GAT_93_ngat), .Y(G537GAT_244_gat) );
AND2XL U_g186 (.A(G506GAT_232_ngat), .B(G317GAT_106_ngat), .Y(G538GAT_245_gat) );
AND2XL U_g187 (.A(G502GAT_234_ngat), .B(G309GAT_107_ngat), .Y(G536GAT_246_gat) );
AND2XL U_g188 (.A(G540GAT_239_gat), .B(G488GAT_184_gat), .Y(G569GAT_247_gat) );
AND2XL U_g189 (.A(G541GAT_238_gat), .B(G489GAT_185_gat), .Y(G573GAT_248_gat) );
AND2XL U_g190 (.A(G542GAT_237_gat), .B(G490GAT_186_gat), .Y(G577GAT_249_gat) );
AND2XL U_g191 (.A(G543GAT_236_gat), .B(G491GAT_187_gat), .Y(G581GAT_250_gat) );
AND2XL U_g192 (.A(G503GAT_203_gat), .B(G536GAT_246_gat), .Y(G553GAT_251_gat) );
AND2XL U_g193 (.A(G505GAT_204_gat), .B(G537GAT_244_gat), .Y(G557GAT_252_gat) );
AND2XL U_g194 (.A(G507GAT_205_gat), .B(G538GAT_245_gat), .Y(G561GAT_253_gat) );
AND2XL U_g195 (.A(G509GAT_206_gat), .B(G539GAT_240_gat), .Y(G565GAT_254_gat) );
BUFX20 U_g196 (.A(G547GAT_235_gat), .Y(G586GAT_255_gat) );
AND2XL U_g197 (.A(G547GAT_235_gat), .B(G544GAT_242_gat), .Y(G587GAT_256_gat) );
BUFX20 U_g198 (.A(G533GAT_241_gat), .Y(G551GAT_257_gat) );
AND2XL U_g199 (.A(G533GAT_241_gat), .B(G530GAT_243_gat), .Y(G552GAT_258_gat) );
BUFX20 U_g200 (.A(G544GAT_242_gat), .Y(G585GAT_259_gat) );
BUFX20 U_g201 (.A(G530GAT_243_gat), .Y(G550GAT_260_gat) );
AND2XL U_g202 (.A(G581GAT_250_gat), .B(G246GAT_53_gat), .Y(G659GAT_261_gat) );
AND2XL U_g203 (.A(G577GAT_249_gat), .B(G246GAT_53_gat), .Y(G650GAT_262_gat) );
AND2XL U_g204 (.A(G573GAT_248_gat), .B(G246GAT_53_gat), .Y(G640GAT_263_gat) );
AND2XL U_g205 (.A(G569GAT_247_gat), .B(G246GAT_53_gat), .Y(G631GAT_264_gat) );
AND2XL U_g206 (.A(G565GAT_254_gat), .B(G246GAT_53_gat), .Y(G624GAT_265_gat) );
AND2XL U_g207 (.A(G561GAT_253_gat), .B(G246GAT_53_gat), .Y(G615GAT_266_gat) );
AND2XL U_g208 (.A(G557GAT_252_gat), .B(G246GAT_53_gat), .Y(G605GAT_267_gat) );
AND2XL U_g209 (.A(G553GAT_251_gat), .B(G246GAT_53_gat), .Y(G596GAT_268_gat) );
AND2XL U_g210 (.A(G586GAT_255_gat), .B(G585GAT_259_gat), .Y(G589GAT_269_gat) );
AND2XL U_g211 (.A(G201GAT_47_ngat), .B(G581GAT_250_ngat), .Y(G654GAT_270_gat) );
AND2XL U_g212 (.A(G201GAT_47_gat), .B(G581GAT_250_gat), .Y(G651GAT_271_gat) );
AND2XL U_g213 (.A(G195GAT_46_ngat), .B(G577GAT_249_ngat), .Y(G644GAT_272_gat) );
AND2XL U_g214 (.A(G195GAT_46_gat), .B(G577GAT_249_gat), .Y(G641GAT_273_gat) );
AND2XL U_g215 (.A(G189GAT_45_ngat), .B(G573GAT_248_ngat), .Y(G635GAT_274_gat) );
AND2XL U_g216 (.A(G189GAT_45_gat), .B(G573GAT_248_gat), .Y(G632GAT_275_gat) );
AND2XL U_g217 (.A(G183GAT_44_ngat), .B(G569GAT_247_ngat), .Y(G628GAT_276_gat) );
AND2XL U_g218 (.A(G183GAT_44_gat), .B(G569GAT_247_gat), .Y(G625GAT_277_gat) );
AND2XL U_g219 (.A(G177GAT_43_ngat), .B(G565GAT_254_ngat), .Y(G619GAT_278_gat) );
AND2XL U_g220 (.A(G177GAT_43_gat), .B(G565GAT_254_gat), .Y(G616GAT_279_gat) );
AND2XL U_g221 (.A(G171GAT_42_ngat), .B(G561GAT_253_ngat), .Y(G609GAT_280_gat) );
AND2XL U_g222 (.A(G171GAT_42_gat), .B(G561GAT_253_gat), .Y(G606GAT_281_gat) );
AND2XL U_g223 (.A(G165GAT_41_ngat), .B(G557GAT_252_ngat), .Y(G600GAT_282_gat) );
AND2XL U_g224 (.A(G165GAT_41_gat), .B(G557GAT_252_gat), .Y(G597GAT_283_gat) );
AND2XL U_g225 (.A(G159GAT_40_ngat), .B(G553GAT_251_ngat), .Y(G593GAT_284_gat) );
AND2XL U_g226 (.A(G159GAT_40_gat), .B(G553GAT_251_gat), .Y(G590GAT_285_gat) );
AND2XL U_g227 (.A(G551GAT_257_gat), .B(G550GAT_260_gat), .Y(G588GAT_286_gat) );
AND4XL U_g228 (.A(G261GAT_57_gat), .B(G654GAT_270_gat), .C(G644GAT_272_gat), .D(G635GAT_274_gat), .Y(G734GAT_287_gat) );
AND3XL U_g229 (.A(G261GAT_57_gat), .B(G654GAT_270_gat), .C(G644GAT_272_gat), .Y(G733GAT_288_gat) );
AND2XL U_g230 (.A(G261GAT_57_gat), .B(G654GAT_270_gat), .Y(G732GAT_289_gat) );
AND2XL U_g231 (.A(G659GAT_261_ngat), .B(G341GAT_61_ngat), .Y(G731GAT_290_gat) );
AND2XL U_g232 (.A(G650GAT_262_ngat), .B(G339GAT_62_ngat), .Y(G721GAT_291_gat) );
AND2XL U_g233 (.A(G640GAT_263_ngat), .B(G337GAT_63_ngat), .Y(G712GAT_292_gat) );
AND2XL U_g234 (.A(G589GAT_269_ngat), .B(G587GAT_256_ngat), .Y(G661GAT_293_gat) );
AND2XL U_g235 (.A(G651GAT_271_gat), .B(G654GAT_270_gat), .Y(G727GAT_294_gat) );
BUFX20 U_g236 (.A(G651GAT_271_gat), .Y(G722GAT_295_gat) );
AND2XL U_g237 (.A(G641GAT_273_gat), .B(G644GAT_272_gat), .Y(G717GAT_296_gat) );
BUFX20 U_g238 (.A(G641GAT_273_gat), .Y(G713GAT_297_gat) );
AND2XL U_g239 (.A(G632GAT_275_gat), .B(G635GAT_274_gat), .Y(G708GAT_298_gat) );
BUFX20 U_g240 (.A(G632GAT_275_gat), .Y(G705GAT_299_gat) );
AND2XL U_g241 (.A(G625GAT_277_gat), .B(G628GAT_276_gat), .Y(G700GAT_300_gat) );
BUFX20 U_g242 (.A(G625GAT_277_gat), .Y(G697GAT_301_gat) );
AND2XL U_g243 (.A(G526GAT_212_ngat), .B(G631GAT_264_ngat), .Y(G704GAT_302_gat) );
AND2XL U_g244 (.A(G616GAT_279_gat), .B(G619GAT_278_gat), .Y(G692GAT_303_gat) );
BUFX20 U_g245 (.A(G616GAT_279_gat), .Y(G687GAT_304_gat) );
AND2XL U_g246 (.A(G525GAT_213_ngat), .B(G624GAT_265_ngat), .Y(G696GAT_305_gat) );
AND2XL U_g247 (.A(G606GAT_281_gat), .B(G609GAT_280_gat), .Y(G682GAT_306_gat) );
BUFX20 U_g248 (.A(G606GAT_281_gat), .Y(G678GAT_307_gat) );
AND2XL U_g249 (.A(G524GAT_214_ngat), .B(G615GAT_266_ngat), .Y(G686GAT_308_gat) );
AND2XL U_g250 (.A(G597GAT_283_gat), .B(G600GAT_282_gat), .Y(G673GAT_309_gat) );
BUFX20 U_g251 (.A(G597GAT_283_gat), .Y(G670GAT_310_gat) );
AND2XL U_g252 (.A(G523GAT_215_ngat), .B(G605GAT_267_ngat), .Y(G677GAT_311_gat) );
AND2XL U_g253 (.A(G590GAT_285_gat), .B(G593GAT_284_gat), .Y(G665GAT_312_gat) );
BUFX20 U_g254 (.A(G590GAT_285_gat), .Y(G662GAT_313_gat) );
AND2XL U_g255 (.A(G522GAT_216_ngat), .B(G596GAT_268_ngat), .Y(G669GAT_314_gat) );
AND2XL U_g256 (.A(G588GAT_286_ngat), .B(G552GAT_258_ngat), .Y(G660GAT_315_gat) );
AND2XL U_g257 (.A(G261GAT_57_gat), .B(G727GAT_294_gat), .Y(G758GAT_316_gat) );
AND2XL U_g258 (.A(G261GAT_57_ngat), .B(G727GAT_294_ngat), .Y(G757GAT_317_gat) );
AND2XL U_g259 (.A(G722GAT_295_gat), .B(G237GAT_52_gat), .Y(G760GAT_318_gat) );
AND2XL U_g260 (.A(G713GAT_297_gat), .B(G237GAT_52_gat), .Y(G755GAT_319_gat) );
AND2XL U_g261 (.A(G705GAT_299_gat), .B(G237GAT_52_gat), .Y(G752GAT_320_gat) );
AND2XL U_g262 (.A(G697GAT_301_gat), .B(G237GAT_52_gat), .Y(G749GAT_321_gat) );
AND2XL U_g263 (.A(G687GAT_304_gat), .B(G237GAT_52_gat), .Y(G746GAT_322_gat) );
AND2XL U_g264 (.A(G678GAT_307_gat), .B(G237GAT_52_gat), .Y(G743GAT_323_gat) );
AND2XL U_g265 (.A(G670GAT_310_gat), .B(G237GAT_52_gat), .Y(G740GAT_324_gat) );
AND2XL U_g266 (.A(G662GAT_313_gat), .B(G237GAT_52_gat), .Y(G737GAT_325_gat) );
AND2XL U_g267 (.A(G727GAT_294_gat), .B(G228GAT_51_gat), .Y(G759GAT_326_gat) );
AND2XL U_g268 (.A(G717GAT_296_gat), .B(G228GAT_51_gat), .Y(G754GAT_327_gat) );
AND2XL U_g269 (.A(G708GAT_298_gat), .B(G228GAT_51_gat), .Y(G751GAT_328_gat) );
AND2XL U_g270 (.A(G700GAT_300_gat), .B(G228GAT_51_gat), .Y(G748GAT_329_gat) );
AND2XL U_g271 (.A(G692GAT_303_gat), .B(G228GAT_51_gat), .Y(G745GAT_330_gat) );
AND2XL U_g272 (.A(G682GAT_306_gat), .B(G228GAT_51_gat), .Y(G742GAT_331_gat) );
AND2XL U_g273 (.A(G673GAT_309_gat), .B(G228GAT_51_gat), .Y(G739GAT_332_gat) );
AND2XL U_g274 (.A(G665GAT_312_gat), .B(G228GAT_51_gat), .Y(G736GAT_333_gat) );
BUFX20 U_g275 (.A(G661GAT_293_gat), .Y(G768GAT_334_gat) );
BUFX20 U_g276 (.A(G722GAT_295_gat), .Y(G756GAT_335_gat) );
AND2XL U_g277 (.A(G722GAT_295_gat), .B(G644GAT_272_gat), .Y(G761GAT_336_gat) );
AND3XL U_g278 (.A(G722GAT_295_gat), .B(G644GAT_272_gat), .C(G635GAT_274_gat), .Y(G763GAT_337_gat) );
BUFX20 U_g279 (.A(G713GAT_297_gat), .Y(G753GAT_338_gat) );
AND2XL U_g280 (.A(G713GAT_297_gat), .B(G635GAT_274_gat), .Y(G762GAT_339_gat) );
BUFX20 U_g281 (.A(G705GAT_299_gat), .Y(G750GAT_340_gat) );
BUFX20 U_g282 (.A(G697GAT_301_gat), .Y(G747GAT_341_gat) );
BUFX20 U_g283 (.A(G687GAT_304_gat), .Y(G744GAT_342_gat) );
AND2XL U_g284 (.A(G687GAT_304_gat), .B(G609GAT_280_gat), .Y(G764GAT_343_gat) );
AND3XL U_g285 (.A(G687GAT_304_gat), .B(G609GAT_280_gat), .C(G600GAT_282_gat), .Y(G766GAT_344_gat) );
BUFX20 U_g286 (.A(G678GAT_307_gat), .Y(G741GAT_345_gat) );
AND2XL U_g287 (.A(G678GAT_307_gat), .B(G600GAT_282_gat), .Y(G765GAT_346_gat) );
BUFX20 U_g288 (.A(G670GAT_310_gat), .Y(G738GAT_347_gat) );
BUFX20 U_g289 (.A(G662GAT_313_gat), .Y(G735GAT_348_gat) );
BUFX20 U_g290 (.A(G660GAT_315_gat), .Y(G767GAT_349_gat) );
AND2XL U_g291 (.A(G758GAT_316_ngat), .B(G757GAT_317_ngat), .Y(G786GAT_350_gat) );
AND4XL U_g292 (.A(G734GAT_287_gat), .B(G763GAT_337_gat), .C(G762GAT_339_gat), .D(G750GAT_340_gat), .Y(G773GAT_351_gat) );
AND3XL U_g293 (.A(G733GAT_288_gat), .B(G761GAT_336_gat), .C(G753GAT_338_gat), .Y(G778GAT_352_gat) );
AND2XL U_g294 (.A(G732GAT_289_gat), .B(G756GAT_335_gat), .Y(G782GAT_353_gat) );
AND2XL U_g295 (.A(G760GAT_318_ngat), .B(G759GAT_326_ngat), .Y(G787GAT_354_gat) );
AND2XL U_g296 (.A(G755GAT_319_ngat), .B(G754GAT_327_ngat), .Y(G785GAT_355_gat) );
AND2XL U_g297 (.A(G752GAT_320_ngat), .B(G751GAT_328_ngat), .Y(G781GAT_356_gat) );
AND2XL U_g298 (.A(G749GAT_321_ngat), .B(G748GAT_329_ngat), .Y(G777GAT_357_gat) );
AND2XL U_g299 (.A(G746GAT_322_ngat), .B(G745GAT_330_ngat), .Y(G772GAT_358_gat) );
AND2XL U_g300 (.A(G743GAT_323_ngat), .B(G742GAT_331_ngat), .Y(G771GAT_359_gat) );
AND2XL U_g301 (.A(G740GAT_324_ngat), .B(G739GAT_332_ngat), .Y(G770GAT_360_gat) );
AND2XL U_g302 (.A(G737GAT_325_ngat), .B(G736GAT_333_ngat), .Y(G769GAT_361_gat) );
AND2XL U_g303 (.A(G786GAT_350_gat), .B(G219GAT_50_gat), .Y(G794GAT_362_gat) );
AND2XL U_g304 (.A(G782GAT_353_ngat), .B(G717GAT_296_ngat), .Y(G792GAT_363_gat) );
AND2XL U_g305 (.A(G782GAT_353_gat), .B(G717GAT_296_gat), .Y(G793GAT_364_gat) );
AND2XL U_g306 (.A(G778GAT_352_ngat), .B(G708GAT_298_ngat), .Y(G790GAT_365_gat) );
AND2XL U_g307 (.A(G778GAT_352_gat), .B(G708GAT_298_gat), .Y(G791GAT_366_gat) );
AND2XL U_g308 (.A(G773GAT_351_ngat), .B(G700GAT_300_ngat), .Y(G788GAT_367_gat) );
AND2XL U_g309 (.A(G773GAT_351_gat), .B(G700GAT_300_gat), .Y(G789GAT_368_gat) );
AND2XL U_g310 (.A(G773GAT_351_gat), .B(G628GAT_276_gat), .Y(G795GAT_369_gat) );
AND2XL U_g311 (.A(G793GAT_364_ngat), .B(G792GAT_363_ngat), .Y(G804GAT_370_gat) );
AND2XL U_g312 (.A(G791GAT_366_ngat), .B(G790GAT_365_ngat), .Y(G803GAT_371_gat) );
AND2XL U_g313 (.A(G789GAT_368_ngat), .B(G788GAT_367_ngat), .Y(G802GAT_372_gat) );
AND2XL U_g314 (.A(G747GAT_341_gat), .B(G795GAT_369_gat), .Y(G796GAT_373_gat) );
AND2XL U_g315 (.A(G794GAT_362_ngat), .B(G340GAT_73_ngat), .Y(G805GAT_374_gat) );
AND2XL U_g316 (.A(G804GAT_370_gat), .B(G219GAT_50_gat), .Y(G810GAT_375_gat) );
AND2XL U_g317 (.A(G803GAT_371_gat), .B(G219GAT_50_gat), .Y(G809GAT_376_gat) );
AND2XL U_g318 (.A(G802GAT_372_gat), .B(G219GAT_50_gat), .Y(G808GAT_377_gat) );
AND4XL U_g319 (.A(G529GAT_209_gat), .B(G731GAT_290_gat), .C(G787GAT_354_gat), .D(G805GAT_374_gat), .Y(G811GAT_378_gat) );
AND2XL U_g320 (.A(G796GAT_373_ngat), .B(G692GAT_303_ngat), .Y(G806GAT_379_gat) );
AND2XL U_g321 (.A(G796GAT_373_gat), .B(G692GAT_303_gat), .Y(G807GAT_380_gat) );
AND2XL U_g322 (.A(G796GAT_373_gat), .B(G619GAT_278_gat), .Y(G812GAT_381_gat) );
AND3XL U_g323 (.A(G796GAT_373_gat), .B(G619GAT_278_gat), .C(G609GAT_280_gat), .Y(G813GAT_382_gat) );
AND4XL U_g324 (.A(G796GAT_373_gat), .B(G619GAT_278_gat), .C(G609GAT_280_gat), .D(G600GAT_282_gat), .Y(G814GAT_383_gat) );
BUFX20 U_g325 (.A(G811GAT_378_gat), .Y(G829GAT_384_gat) );
AND2XL U_g326 (.A(G807GAT_380_ngat), .B(G806GAT_379_ngat), .Y(G825GAT_385_gat) );
AND2XL U_g327 (.A(G812GAT_381_gat), .B(G744GAT_342_gat), .Y(G822GAT_386_gat) );
AND3XL U_g328 (.A(G813GAT_382_gat), .B(G764GAT_343_gat), .C(G741GAT_345_gat), .Y(G819GAT_387_gat) );
AND4XL U_g329 (.A(G814GAT_383_gat), .B(G766GAT_344_gat), .C(G765GAT_346_gat), .D(G738GAT_347_gat), .Y(G815GAT_388_gat) );
AND2XL U_g330 (.A(G810GAT_375_ngat), .B(G338GAT_76_ngat), .Y(G828GAT_389_gat) );
AND2XL U_g331 (.A(G809GAT_376_ngat), .B(G336GAT_77_ngat), .Y(G827GAT_390_gat) );
AND2XL U_g332 (.A(G808GAT_377_ngat), .B(G335GAT_80_ngat), .Y(G826GAT_391_gat) );
AND2XL U_g333 (.A(G825GAT_385_gat), .B(G219GAT_50_gat), .Y(G836GAT_392_gat) );
BUFX20 U_g334 (.A(G829GAT_384_gat), .Y(G840GAT_393_gat) );
AND4XL U_g335 (.A(G528GAT_210_gat), .B(G721GAT_291_gat), .C(G785GAT_355_gat), .D(G828GAT_389_gat), .Y(G839GAT_394_gat) );
AND4XL U_g336 (.A(G527GAT_211_gat), .B(G712GAT_292_gat), .C(G781GAT_356_gat), .D(G827GAT_390_gat), .Y(G838GAT_395_gat) );
AND3XL U_g337 (.A(G704GAT_302_gat), .B(G777GAT_357_gat), .C(G826GAT_391_gat), .Y(G837GAT_396_gat) );
AND2XL U_g338 (.A(G822GAT_386_ngat), .B(G682GAT_306_ngat), .Y(G834GAT_397_gat) );
AND2XL U_g339 (.A(G822GAT_386_gat), .B(G682GAT_306_gat), .Y(G835GAT_398_gat) );
AND2XL U_g340 (.A(G819GAT_387_ngat), .B(G673GAT_309_ngat), .Y(G832GAT_399_gat) );
AND2XL U_g341 (.A(G819GAT_387_gat), .B(G673GAT_309_gat), .Y(G833GAT_400_gat) );
AND2XL U_g342 (.A(G815GAT_388_ngat), .B(G665GAT_312_ngat), .Y(G830GAT_401_gat) );
AND2XL U_g343 (.A(G815GAT_388_gat), .B(G665GAT_312_gat), .Y(G831GAT_402_gat) );
AND2XL U_g344 (.A(G593GAT_284_gat), .B(G815GAT_388_gat), .Y(G841GAT_403_gat) );
BUFX20 U_g345 (.A(G840GAT_393_gat), .Y(G850GAT_404_gat) );
BUFX20 U_g346 (.A(G839GAT_394_gat), .Y(G848GAT_405_gat) );
BUFX20 U_g347 (.A(G838GAT_395_gat), .Y(G847GAT_406_gat) );
BUFX20 U_g348 (.A(G837GAT_396_gat), .Y(G846GAT_407_gat) );
AND2XL U_g349 (.A(G835GAT_398_ngat), .B(G834GAT_397_ngat), .Y(G844GAT_408_gat) );
AND2XL U_g350 (.A(G833GAT_400_ngat), .B(G832GAT_399_ngat), .Y(G843GAT_409_gat) );
AND2XL U_g351 (.A(G831GAT_402_ngat), .B(G830GAT_401_ngat), .Y(G842GAT_410_gat) );
AND2XL U_g352 (.A(G841GAT_403_gat), .B(G735GAT_348_gat), .Y(G849GAT_411_gat) );
AND2XL U_g353 (.A(G836GAT_392_ngat), .B(G334GAT_81_ngat), .Y(G845GAT_412_gat) );
AND2XL U_g354 (.A(G844GAT_408_gat), .B(G219GAT_50_gat), .Y(G853GAT_413_gat) );
AND2XL U_g355 (.A(G843GAT_409_gat), .B(G219GAT_50_gat), .Y(G852GAT_414_gat) );
AND2XL U_g356 (.A(G842GAT_410_gat), .B(G219GAT_50_gat), .Y(G851GAT_415_gat) );
BUFX20 U_g357 (.A(G848GAT_405_gat), .Y(G857GAT_416_gat) );
BUFX20 U_g358 (.A(G847GAT_406_gat), .Y(G856GAT_417_gat) );
BUFX20 U_g359 (.A(G846GAT_407_gat), .Y(G855GAT_418_gat) );
AND3XL U_g360 (.A(G696GAT_305_gat), .B(G772GAT_358_gat), .C(G845GAT_412_gat), .Y(G854GAT_419_gat) );
BUFX20 U_g361 (.A(G849GAT_411_gat), .Y(G858GAT_420_gat) );
AND2XL U_g362 (.A(G851GAT_415_ngat), .B(G417GAT_142_ngat), .Y(G859GAT_421_gat) );
BUFX20 U_g363 (.A(G857GAT_416_gat), .Y(G865GAT_422_gat) );
BUFX20 U_g364 (.A(G856GAT_417_gat), .Y(G864GAT_423_gat) );
BUFX20 U_g365 (.A(G855GAT_418_gat), .Y(G863GAT_424_gat) );
BUFX20 U_g366 (.A(G854GAT_419_gat), .Y(G862GAT_425_gat) );
BUFX20 U_g367 (.A(G858GAT_420_gat), .Y(G866GAT_426_gat) );
AND2XL U_g368 (.A(G853GAT_413_ngat), .B(G333GAT_84_ngat), .Y(G861GAT_427_gat) );
AND2XL U_g369 (.A(G852GAT_414_ngat), .B(G332GAT_85_ngat), .Y(G860GAT_428_gat) );
BUFX20 U_g370 (.A(G862GAT_425_gat), .Y(G870GAT_429_gat) );
AND3XL U_g371 (.A(G686GAT_308_gat), .B(G771GAT_359_gat), .C(G861GAT_427_gat), .Y(G869GAT_430_gat) );
AND3XL U_g372 (.A(G677GAT_311_gat), .B(G770GAT_360_gat), .C(G860GAT_428_gat), .Y(G868GAT_431_gat) );
AND3XL U_g373 (.A(G669GAT_314_gat), .B(G769GAT_361_gat), .C(G859GAT_421_gat), .Y(G867GAT_432_gat) );
BUFX20 U_g374 (.A(G870GAT_429_gat), .Y(G874GAT_433_gat) );
BUFX20 U_g375 (.A(G869GAT_430_gat), .Y(G873GAT_434_gat) );
BUFX20 U_g376 (.A(G868GAT_431_gat), .Y(G872GAT_435_gat) );
BUFX20 U_g377 (.A(G867GAT_432_gat), .Y(G871GAT_436_gat) );
BUFX20 U_g378 (.A(G873GAT_434_gat), .Y(G877GAT_437_gat) );
BUFX20 U_g379 (.A(G872GAT_435_gat), .Y(G876GAT_438_gat) );
BUFX20 U_g380 (.A(G871GAT_436_gat), .Y(G875GAT_439_gat) );
BUFX20 U_g381 (.A(G877GAT_437_gat), .Y(G880GAT_440_gat) );
BUFX20 U_g382 (.A(G876GAT_438_gat), .Y(G879GAT_441_gat) );
BUFX20 U_g383 (.A(G875GAT_439_gat), .Y(G878GAT_442_gat) );
INVXL U_g384 (.A(G195GAT_46_gat), .Y(G195GAT_46_ngat) );
INVXL U_g385 (.A(G201GAT_47_gat), .Y(G201GAT_47_ngat) );
INVXL U_g386 (.A(G183GAT_44_gat), .Y(G183GAT_44_ngat) );
INVXL U_g387 (.A(G189GAT_45_gat), .Y(G189GAT_45_ngat) );
INVXL U_g388 (.A(G171GAT_42_gat), .Y(G171GAT_42_ngat) );
INVXL U_g389 (.A(G177GAT_43_gat), .Y(G177GAT_43_ngat) );
INVXL U_g390 (.A(G159GAT_40_gat), .Y(G159GAT_40_ngat) );
INVXL U_g391 (.A(G165GAT_41_gat), .Y(G165GAT_41_ngat) );
INVXL U_g392 (.A(G121GAT_29_gat), .Y(G121GAT_29_ngat) );
INVXL U_g393 (.A(G126GAT_30_gat), .Y(G126GAT_30_ngat) );
INVXL U_g394 (.A(G111GAT_27_gat), .Y(G111GAT_27_ngat) );
INVXL U_g395 (.A(G116GAT_28_gat), .Y(G116GAT_28_ngat) );
INVXL U_g396 (.A(G101GAT_25_gat), .Y(G101GAT_25_ngat) );
INVXL U_g397 (.A(G106GAT_26_gat), .Y(G106GAT_26_ngat) );
INVXL U_g398 (.A(G91GAT_23_gat), .Y(G91GAT_23_ngat) );
INVXL U_g399 (.A(G96GAT_24_gat), .Y(G96GAT_24_ngat) );
INVXL U_g400 (.A(G87GAT_19_gat), .Y(G87GAT_19_ngat) );
INVXL U_g401 (.A(G88GAT_20_gat), .Y(G88GAT_20_ngat) );
INVXL U_g402 (.A(G17GAT_3_gat), .Y(G17GAT_3_ngat) );
INVXL U_g403 (.A(G42GAT_7_gat), .Y(G42GAT_7_ngat) );
INVXL U_g404 (.A(G280GAT_108_gat), .Y(G280GAT_108_ngat) );
INVXL U_g405 (.A(G286GAT_92_gat), .Y(G286GAT_92_ngat) );
INVXL U_g406 (.A(G284GAT_95_gat), .Y(G284GAT_95_ngat) );
INVXL U_g407 (.A(G285GAT_102_gat), .Y(G285GAT_102_ngat) );
INVXL U_g408 (.A(G270GAT_111_gat), .Y(G270GAT_111_ngat) );
INVXL U_g409 (.A(G273GAT_103_gat), .Y(G273GAT_103_ngat) );
INVXL U_g410 (.A(G322GAT_105_gat), .Y(G322GAT_105_ngat) );
INVXL U_g411 (.A(G323GAT_104_gat), .Y(G323GAT_104_ngat) );
INVXL U_g412 (.A(G343GAT_135_gat), .Y(G343GAT_135_ngat) );
INVXL U_g413 (.A(G369GAT_113_gat), .Y(G369GAT_113_ngat) );
INVXL U_g414 (.A(G437GAT_177_gat), .Y(G437GAT_177_ngat) );
INVXL U_g415 (.A(G416GAT_144_gat), .Y(G416GAT_144_ngat) );
INVXL U_g416 (.A(G445GAT_169_gat), .Y(G445GAT_169_ngat) );
INVXL U_g417 (.A(G413GAT_147_gat), .Y(G413GAT_147_ngat) );
INVXL U_g418 (.A(G444GAT_170_gat), .Y(G444GAT_170_ngat) );
INVXL U_g419 (.A(G409GAT_150_gat), .Y(G409GAT_150_ngat) );
INVXL U_g420 (.A(G426GAT_171_gat), .Y(G426GAT_171_ngat) );
INVXL U_g421 (.A(G406GAT_153_gat), .Y(G406GAT_153_ngat) );
INVXL U_g422 (.A(G425GAT_172_gat), .Y(G425GAT_172_ngat) );
INVXL U_g423 (.A(G475GAT_197_gat), .Y(G475GAT_197_ngat) );
INVXL U_g424 (.A(G476GAT_188_gat), .Y(G476GAT_188_ngat) );
INVXL U_g425 (.A(G477GAT_196_gat), .Y(G477GAT_196_ngat) );
INVXL U_g426 (.A(G478GAT_189_gat), .Y(G478GAT_189_ngat) );
INVXL U_g427 (.A(G479GAT_195_gat), .Y(G479GAT_195_ngat) );
INVXL U_g428 (.A(G480GAT_190_gat), .Y(G480GAT_190_ngat) );
INVXL U_g429 (.A(G481GAT_194_gat), .Y(G481GAT_194_ngat) );
INVXL U_g430 (.A(G482GAT_191_gat), .Y(G482GAT_191_ngat) );
INVXL U_g431 (.A(G495GAT_192_gat), .Y(G495GAT_192_ngat) );
INVXL U_g432 (.A(G207GAT_48_gat), .Y(G207GAT_48_ngat) );
INVXL U_g433 (.A(G463GAT_198_gat), .Y(G463GAT_198_ngat) );
INVXL U_g434 (.A(G135GAT_32_gat), .Y(G135GAT_32_ngat) );
INVXL U_g435 (.A(G130GAT_31_gat), .Y(G130GAT_31_ngat) );
INVXL U_g436 (.A(G492GAT_193_gat), .Y(G492GAT_193_ngat) );
INVXL U_g437 (.A(G460GAT_199_gat), .Y(G460GAT_199_ngat) );
INVXL U_g438 (.A(G516GAT_217_gat), .Y(G516GAT_217_ngat) );
INVXL U_g439 (.A(G517GAT_227_gat), .Y(G517GAT_227_ngat) );
INVXL U_g440 (.A(G514GAT_218_gat), .Y(G514GAT_218_ngat) );
INVXL U_g441 (.A(G515GAT_228_gat), .Y(G515GAT_228_ngat) );
INVXL U_g442 (.A(G512GAT_219_gat), .Y(G512GAT_219_ngat) );
INVXL U_g443 (.A(G513GAT_229_gat), .Y(G513GAT_229_ngat) );
INVXL U_g444 (.A(G510GAT_220_gat), .Y(G510GAT_220_ngat) );
INVXL U_g445 (.A(G511GAT_230_gat), .Y(G511GAT_230_ngat) );
INVXL U_g446 (.A(G318GAT_72_gat), .Y(G318GAT_72_ngat) );
INVXL U_g447 (.A(G508GAT_231_gat), .Y(G508GAT_231_ngat) );
INVXL U_g448 (.A(G316GAT_93_gat), .Y(G316GAT_93_ngat) );
INVXL U_g449 (.A(G504GAT_233_gat), .Y(G504GAT_233_ngat) );
INVXL U_g450 (.A(G317GAT_106_gat), .Y(G317GAT_106_ngat) );
INVXL U_g451 (.A(G506GAT_232_gat), .Y(G506GAT_232_ngat) );
INVXL U_g452 (.A(G309GAT_107_gat), .Y(G309GAT_107_ngat) );
INVXL U_g453 (.A(G502GAT_234_gat), .Y(G502GAT_234_ngat) );
INVXL U_g454 (.A(G581GAT_250_gat), .Y(G581GAT_250_ngat) );
INVXL U_g455 (.A(G577GAT_249_gat), .Y(G577GAT_249_ngat) );
INVXL U_g456 (.A(G573GAT_248_gat), .Y(G573GAT_248_ngat) );
INVXL U_g457 (.A(G569GAT_247_gat), .Y(G569GAT_247_ngat) );
INVXL U_g458 (.A(G565GAT_254_gat), .Y(G565GAT_254_ngat) );
INVXL U_g459 (.A(G561GAT_253_gat), .Y(G561GAT_253_ngat) );
INVXL U_g460 (.A(G557GAT_252_gat), .Y(G557GAT_252_ngat) );
INVXL U_g461 (.A(G553GAT_251_gat), .Y(G553GAT_251_ngat) );
INVXL U_g462 (.A(G341GAT_61_gat), .Y(G341GAT_61_ngat) );
INVXL U_g463 (.A(G659GAT_261_gat), .Y(G659GAT_261_ngat) );
INVXL U_g464 (.A(G339GAT_62_gat), .Y(G339GAT_62_ngat) );
INVXL U_g465 (.A(G650GAT_262_gat), .Y(G650GAT_262_ngat) );
INVXL U_g466 (.A(G337GAT_63_gat), .Y(G337GAT_63_ngat) );
INVXL U_g467 (.A(G640GAT_263_gat), .Y(G640GAT_263_ngat) );
INVXL U_g468 (.A(G587GAT_256_gat), .Y(G587GAT_256_ngat) );
INVXL U_g469 (.A(G589GAT_269_gat), .Y(G589GAT_269_ngat) );
INVXL U_g470 (.A(G631GAT_264_gat), .Y(G631GAT_264_ngat) );
INVXL U_g471 (.A(G526GAT_212_gat), .Y(G526GAT_212_ngat) );
INVXL U_g472 (.A(G624GAT_265_gat), .Y(G624GAT_265_ngat) );
INVXL U_g473 (.A(G525GAT_213_gat), .Y(G525GAT_213_ngat) );
INVXL U_g474 (.A(G615GAT_266_gat), .Y(G615GAT_266_ngat) );
INVXL U_g475 (.A(G524GAT_214_gat), .Y(G524GAT_214_ngat) );
INVXL U_g476 (.A(G605GAT_267_gat), .Y(G605GAT_267_ngat) );
INVXL U_g477 (.A(G523GAT_215_gat), .Y(G523GAT_215_ngat) );
INVXL U_g478 (.A(G596GAT_268_gat), .Y(G596GAT_268_ngat) );
INVXL U_g479 (.A(G522GAT_216_gat), .Y(G522GAT_216_ngat) );
INVXL U_g480 (.A(G552GAT_258_gat), .Y(G552GAT_258_ngat) );
INVXL U_g481 (.A(G588GAT_286_gat), .Y(G588GAT_286_ngat) );
INVXL U_g482 (.A(G727GAT_294_gat), .Y(G727GAT_294_ngat) );
INVXL U_g483 (.A(G261GAT_57_gat), .Y(G261GAT_57_ngat) );
INVXL U_g484 (.A(G757GAT_317_gat), .Y(G757GAT_317_ngat) );
INVXL U_g485 (.A(G758GAT_316_gat), .Y(G758GAT_316_ngat) );
INVXL U_g486 (.A(G759GAT_326_gat), .Y(G759GAT_326_ngat) );
INVXL U_g487 (.A(G760GAT_318_gat), .Y(G760GAT_318_ngat) );
INVXL U_g488 (.A(G754GAT_327_gat), .Y(G754GAT_327_ngat) );
INVXL U_g489 (.A(G755GAT_319_gat), .Y(G755GAT_319_ngat) );
INVXL U_g490 (.A(G751GAT_328_gat), .Y(G751GAT_328_ngat) );
INVXL U_g491 (.A(G752GAT_320_gat), .Y(G752GAT_320_ngat) );
INVXL U_g492 (.A(G748GAT_329_gat), .Y(G748GAT_329_ngat) );
INVXL U_g493 (.A(G749GAT_321_gat), .Y(G749GAT_321_ngat) );
INVXL U_g494 (.A(G745GAT_330_gat), .Y(G745GAT_330_ngat) );
INVXL U_g495 (.A(G746GAT_322_gat), .Y(G746GAT_322_ngat) );
INVXL U_g496 (.A(G742GAT_331_gat), .Y(G742GAT_331_ngat) );
INVXL U_g497 (.A(G743GAT_323_gat), .Y(G743GAT_323_ngat) );
INVXL U_g498 (.A(G739GAT_332_gat), .Y(G739GAT_332_ngat) );
INVXL U_g499 (.A(G740GAT_324_gat), .Y(G740GAT_324_ngat) );
INVXL U_g500 (.A(G736GAT_333_gat), .Y(G736GAT_333_ngat) );
INVXL U_g501 (.A(G737GAT_325_gat), .Y(G737GAT_325_ngat) );
INVXL U_g502 (.A(G717GAT_296_gat), .Y(G717GAT_296_ngat) );
INVXL U_g503 (.A(G782GAT_353_gat), .Y(G782GAT_353_ngat) );
INVXL U_g504 (.A(G708GAT_298_gat), .Y(G708GAT_298_ngat) );
INVXL U_g505 (.A(G778GAT_352_gat), .Y(G778GAT_352_ngat) );
INVXL U_g506 (.A(G700GAT_300_gat), .Y(G700GAT_300_ngat) );
INVXL U_g507 (.A(G773GAT_351_gat), .Y(G773GAT_351_ngat) );
INVXL U_g508 (.A(G792GAT_363_gat), .Y(G792GAT_363_ngat) );
INVXL U_g509 (.A(G793GAT_364_gat), .Y(G793GAT_364_ngat) );
INVXL U_g510 (.A(G790GAT_365_gat), .Y(G790GAT_365_ngat) );
INVXL U_g511 (.A(G791GAT_366_gat), .Y(G791GAT_366_ngat) );
INVXL U_g512 (.A(G788GAT_367_gat), .Y(G788GAT_367_ngat) );
INVXL U_g513 (.A(G789GAT_368_gat), .Y(G789GAT_368_ngat) );
INVXL U_g514 (.A(G340GAT_73_gat), .Y(G340GAT_73_ngat) );
INVXL U_g515 (.A(G794GAT_362_gat), .Y(G794GAT_362_ngat) );
INVXL U_g516 (.A(G692GAT_303_gat), .Y(G692GAT_303_ngat) );
INVXL U_g517 (.A(G796GAT_373_gat), .Y(G796GAT_373_ngat) );
INVXL U_g518 (.A(G806GAT_379_gat), .Y(G806GAT_379_ngat) );
INVXL U_g519 (.A(G807GAT_380_gat), .Y(G807GAT_380_ngat) );
INVXL U_g520 (.A(G338GAT_76_gat), .Y(G338GAT_76_ngat) );
INVXL U_g521 (.A(G810GAT_375_gat), .Y(G810GAT_375_ngat) );
INVXL U_g522 (.A(G336GAT_77_gat), .Y(G336GAT_77_ngat) );
INVXL U_g523 (.A(G809GAT_376_gat), .Y(G809GAT_376_ngat) );
INVXL U_g524 (.A(G335GAT_80_gat), .Y(G335GAT_80_ngat) );
INVXL U_g525 (.A(G808GAT_377_gat), .Y(G808GAT_377_ngat) );
INVXL U_g526 (.A(G682GAT_306_gat), .Y(G682GAT_306_ngat) );
INVXL U_g527 (.A(G822GAT_386_gat), .Y(G822GAT_386_ngat) );
INVXL U_g528 (.A(G673GAT_309_gat), .Y(G673GAT_309_ngat) );
INVXL U_g529 (.A(G819GAT_387_gat), .Y(G819GAT_387_ngat) );
INVXL U_g530 (.A(G665GAT_312_gat), .Y(G665GAT_312_ngat) );
INVXL U_g531 (.A(G815GAT_388_gat), .Y(G815GAT_388_ngat) );
INVXL U_g532 (.A(G834GAT_397_gat), .Y(G834GAT_397_ngat) );
INVXL U_g533 (.A(G835GAT_398_gat), .Y(G835GAT_398_ngat) );
INVXL U_g534 (.A(G832GAT_399_gat), .Y(G832GAT_399_ngat) );
INVXL U_g535 (.A(G833GAT_400_gat), .Y(G833GAT_400_ngat) );
INVXL U_g536 (.A(G830GAT_401_gat), .Y(G830GAT_401_ngat) );
INVXL U_g537 (.A(G831GAT_402_gat), .Y(G831GAT_402_ngat) );
INVXL U_g538 (.A(G334GAT_81_gat), .Y(G334GAT_81_ngat) );
INVXL U_g539 (.A(G836GAT_392_gat), .Y(G836GAT_392_ngat) );
INVXL U_g540 (.A(G417GAT_142_gat), .Y(G417GAT_142_ngat) );
INVXL U_g541 (.A(G851GAT_415_gat), .Y(G851GAT_415_ngat) );
INVXL U_g542 (.A(G333GAT_84_gat), .Y(G333GAT_84_ngat) );
INVXL U_g543 (.A(G853GAT_413_gat), .Y(G853GAT_413_ngat) );
INVXL U_g544 (.A(G332GAT_85_gat), .Y(G332GAT_85_ngat) );
INVXL U_g545 (.A(G852GAT_414_gat), .Y(G852GAT_414_ngat) );

endmodule
