module C2670 ( G1_0_gat, G2_1_gat, G3_2_gat, G4_3_gat, G5_4_gat, G6_5_gat, G7_6_gat, G8_7_gat, G11_8_gat, G14_9_gat, G15_10_gat, G16_11_gat, G19_12_gat, G20_13_gat, G21_14_gat, G22_15_gat, G23_16_gat, G24_17_gat, G25_18_gat, G26_19_gat, G27_20_gat, G28_21_gat, G29_22_gat, G32_23_gat, G33_24_gat, G34_25_gat, G35_26_gat, G36_27_gat, G37_28_gat, G40_29_gat, G43_30_gat, G44_31_gat, G47_32_gat, G48_33_gat, G49_34_gat, G50_35_gat, G51_36_gat, G52_37_gat, G53_38_gat, G54_39_gat, G55_40_gat, G56_41_gat, G57_42_gat, G60_43_gat, G61_44_gat, G62_45_gat, G63_46_gat, G64_47_gat, G65_48_gat, G66_49_gat, G67_50_gat, G68_51_gat, G69_52_gat, G72_53_gat, G73_54_gat, G74_55_gat, G75_56_gat, G76_57_gat, G77_58_gat, G78_59_gat, G79_60_gat, G80_61_gat, G81_62_gat, G82_63_gat, G85_64_gat, G86_65_gat, G87_66_gat, G88_67_gat, G89_68_gat, G90_69_gat, G91_70_gat, G92_71_gat, G93_72_gat, G94_73_gat, G95_74_gat, G96_75_gat, G99_76_gat, G100_77_gat, G101_78_gat, G102_79_gat, G103_80_gat, G104_81_gat, G105_82_gat, G106_83_gat, G107_84_gat, G108_85_gat, G111_86_gat, G112_87_gat, G113_88_gat, G114_89_gat, G115_90_gat, G116_91_gat, G117_92_gat, G118_93_gat, G119_94_gat, G120_95_gat, G123_96_gat, G124_97_gat, G125_98_gat, G126_99_gat, G127_100_gat, G128_101_gat, G129_102_gat, G130_103_gat, G131_104_gat, G132_105_gat, G135_106_gat, G136_107_gat, G137_108_gat, G138_109_gat, G139_110_gat, G140_111_gat, G141_112_gat, G142_113_gat, GIN_169_114_gat, GIN_174_115_gat, GIN_177_116_gat, GIN_178_117_gat, GIN_179_118_gat, GIN_180_119_gat, GIN_181_120_gat, GIN_182_121_gat, GIN_183_122_gat, GIN_184_123_gat, GIN_185_124_gat, GIN_186_125_gat, GIN_189_126_gat, GIN_190_127_gat, GIN_191_128_gat, GIN_192_129_gat, GIN_193_130_gat, GIN_194_131_gat, GIN_195_132_gat, GIN_196_133_gat, GIN_197_134_gat, GIN_198_135_gat, GIN_199_136_gat, GIN_200_137_gat, GIN_201_138_gat, GIN_202_139_gat, GIN_203_140_gat, GIN_204_141_gat, GIN_205_142_gat, GIN_206_143_gat, GIN_207_144_gat, GIN_208_145_gat, GIN_209_146_gat, GIN_210_147_gat, GIN_211_148_gat, GIN_212_149_gat, GIN_213_150_gat, GIN_214_151_gat, GIN_215_152_gat, GIN_239_153_gat, GIN_240_154_gat, GIN_241_155_gat, GIN_242_156_gat, GIN_243_157_gat, GIN_244_158_gat, GIN_245_159_gat, GIN_246_160_gat, GIN_247_161_gat, GIN_248_162_gat, GIN_249_163_gat, GIN_250_164_gat, GIN_251_165_gat, GIN_252_166_gat, GIN_253_167_gat, GIN_254_168_gat, GIN_255_169_gat, GIN_256_170_gat, GIN_257_171_gat, GIN_262_172_gat, GIN_263_173_gat, GIN_264_174_gat, GIN_265_175_gat, GIN_266_176_gat, GIN_267_177_gat, GIN_268_178_gat, GIN_269_179_gat, GIN_270_180_gat, GIN_271_181_gat, GIN_272_182_gat, GIN_273_183_gat, GIN_274_184_gat, GIN_275_185_gat, GIN_276_186_gat, GIN_277_187_gat, GIN_278_188_gat, GIN_279_189_gat, G452_190_gat, G483_191_gat, G543_192_gat, G559_193_gat, G567_194_gat, G651_195_gat, G661_196_gat, G860_197_gat, G868_198_gat, G1083_199_gat, G1341_200_gat, G1348_201_gat, G1384_202_gat, G1956_203_gat, G1961_204_gat, G1966_205_gat, G1971_206_gat, G1976_207_gat, G1981_208_gat, G1986_209_gat, G1991_210_gat, G1996_211_gat, G2066_212_gat, G2067_213_gat, G2072_214_gat, G2078_215_gat, G2084_216_gat, G2090_217_gat, G2096_218_gat, G2100_219_gat, G2104_220_gat, G2105_221_gat, G2106_222_gat, G2427_223_gat, G2430_224_gat, G2435_225_gat, G2438_226_gat, G2443_227_gat, G2446_228_gat, G2451_229_gat, G2454_230_gat, G2474_231_gat, G2678_232_gat, G169_114_gat, G174_115_gat, G177_116_gat, G178_117_gat, G179_118_gat, G180_119_gat, G181_120_gat, G182_121_gat, G183_122_gat, G184_123_gat, G185_124_gat, G186_125_gat, G189_126_gat, G190_127_gat, G191_128_gat, G192_129_gat, G193_130_gat, G194_131_gat, G195_132_gat, G196_133_gat, G197_134_gat, G198_135_gat, G199_136_gat, G200_137_gat, G201_138_gat, G202_139_gat, G203_140_gat, G204_141_gat, G205_142_gat, G206_143_gat, G207_144_gat, G208_145_gat, G209_146_gat, G210_147_gat, G211_148_gat, G212_149_gat, G213_150_gat, G214_151_gat, G215_152_gat, G239_153_gat, G240_154_gat, G241_155_gat, G242_156_gat, G243_157_gat, G244_158_gat, G245_159_gat, G246_160_gat, G247_161_gat, G248_162_gat, G249_163_gat, G250_164_gat, G251_165_gat, G252_166_gat, G253_167_gat, G254_168_gat, G255_169_gat, G256_170_gat, G257_171_gat, G262_172_gat, G263_173_gat, G264_174_gat, G265_175_gat, G266_176_gat, G267_177_gat, G268_178_gat, G269_179_gat, G270_180_gat, G271_181_gat, G272_182_gat, G273_183_gat, G274_184_gat, G275_185_gat, G276_186_gat, G277_187_gat, G278_188_gat, G279_189_gat, G350_301_gat, G335_299_gat, G409_298_gat, G369_289_gat, G367_288_gat, G411_264_gat, G337_263_gat, G384_262_gat, G218_311_gat, G219_302_gat, G220_306_gat, G221_305_gat, G235_307_gat, G236_303_gat, G237_309_gat, G238_304_gat, G158_349_gat, G259_414_gat, G391_379_gat, G173_389_gat, G223_413_gat, G234_376_gat, G217_423_gat, G325_507_gat, G261_506_gat, G319_656_gat, G160_609_gat, G162_612_gat, G164_607_gat, G166_625_gat, G168_623_gat, G171_621_gat, G153_671_gat, G176_803_gat, G188_761_gat, G299_692_gat, G301_694_gat, G286_696_gat, G303_698_gat, G288_700_gat, G305_702_gat, G290_704_gat, G284_847_gat, G321_848_gat, G297_849_gat, G280_850_gat, G148_851_gat, G282_922_gat, G323_923_gat, G156_1046_gat, G401_1276_gat, G227_1179_gat, G229_1180_gat, G311_1278_gat, G150_1277_gat, G145_1358_gat, G395_1392_gat, G295_1400_gat, G331_1401_gat, G397_1406_gat, G329_1414_gat, G231_1422_gat, G308_1425_gat, G225_1424_gat);

input G1_0_gat;
input G2_1_gat;
input G3_2_gat;
input G4_3_gat;
input G5_4_gat;
input G6_5_gat;
input G7_6_gat;
input G8_7_gat;
input G11_8_gat;
input G14_9_gat;
input G15_10_gat;
input G16_11_gat;
input G19_12_gat;
input G20_13_gat;
input G21_14_gat;
input G22_15_gat;
input G23_16_gat;
input G24_17_gat;
input G25_18_gat;
input G26_19_gat;
input G27_20_gat;
input G28_21_gat;
input G29_22_gat;
input G32_23_gat;
input G33_24_gat;
input G34_25_gat;
input G35_26_gat;
input G36_27_gat;
input G37_28_gat;
input G40_29_gat;
input G43_30_gat;
input G44_31_gat;
input G47_32_gat;
input G48_33_gat;
input G49_34_gat;
input G50_35_gat;
input G51_36_gat;
input G52_37_gat;
input G53_38_gat;
input G54_39_gat;
input G55_40_gat;
input G56_41_gat;
input G57_42_gat;
input G60_43_gat;
input G61_44_gat;
input G62_45_gat;
input G63_46_gat;
input G64_47_gat;
input G65_48_gat;
input G66_49_gat;
input G67_50_gat;
input G68_51_gat;
input G69_52_gat;
input G72_53_gat;
input G73_54_gat;
input G74_55_gat;
input G75_56_gat;
input G76_57_gat;
input G77_58_gat;
input G78_59_gat;
input G79_60_gat;
input G80_61_gat;
input G81_62_gat;
input G82_63_gat;
input G85_64_gat;
input G86_65_gat;
input G87_66_gat;
input G88_67_gat;
input G89_68_gat;
input G90_69_gat;
input G91_70_gat;
input G92_71_gat;
input G93_72_gat;
input G94_73_gat;
input G95_74_gat;
input G96_75_gat;
input G99_76_gat;
input G100_77_gat;
input G101_78_gat;
input G102_79_gat;
input G103_80_gat;
input G104_81_gat;
input G105_82_gat;
input G106_83_gat;
input G107_84_gat;
input G108_85_gat;
input G111_86_gat;
input G112_87_gat;
input G113_88_gat;
input G114_89_gat;
input G115_90_gat;
input G116_91_gat;
input G117_92_gat;
input G118_93_gat;
input G119_94_gat;
input G120_95_gat;
input G123_96_gat;
input G124_97_gat;
input G125_98_gat;
input G126_99_gat;
input G127_100_gat;
input G128_101_gat;
input G129_102_gat;
input G130_103_gat;
input G131_104_gat;
input G132_105_gat;
input G135_106_gat;
input G136_107_gat;
input G137_108_gat;
input G138_109_gat;
input G139_110_gat;
input G140_111_gat;
input G141_112_gat;
input G142_113_gat;
input GIN_169_114_gat;
input GIN_174_115_gat;
input GIN_177_116_gat;
input GIN_178_117_gat;
input GIN_179_118_gat;
input GIN_180_119_gat;
input GIN_181_120_gat;
input GIN_182_121_gat;
input GIN_183_122_gat;
input GIN_184_123_gat;
input GIN_185_124_gat;
input GIN_186_125_gat;
input GIN_189_126_gat;
input GIN_190_127_gat;
input GIN_191_128_gat;
input GIN_192_129_gat;
input GIN_193_130_gat;
input GIN_194_131_gat;
input GIN_195_132_gat;
input GIN_196_133_gat;
input GIN_197_134_gat;
input GIN_198_135_gat;
input GIN_199_136_gat;
input GIN_200_137_gat;
input GIN_201_138_gat;
input GIN_202_139_gat;
input GIN_203_140_gat;
input GIN_204_141_gat;
input GIN_205_142_gat;
input GIN_206_143_gat;
input GIN_207_144_gat;
input GIN_208_145_gat;
input GIN_209_146_gat;
input GIN_210_147_gat;
input GIN_211_148_gat;
input GIN_212_149_gat;
input GIN_213_150_gat;
input GIN_214_151_gat;
input GIN_215_152_gat;
input GIN_239_153_gat;
input GIN_240_154_gat;
input GIN_241_155_gat;
input GIN_242_156_gat;
input GIN_243_157_gat;
input GIN_244_158_gat;
input GIN_245_159_gat;
input GIN_246_160_gat;
input GIN_247_161_gat;
input GIN_248_162_gat;
input GIN_249_163_gat;
input GIN_250_164_gat;
input GIN_251_165_gat;
input GIN_252_166_gat;
input GIN_253_167_gat;
input GIN_254_168_gat;
input GIN_255_169_gat;
input GIN_256_170_gat;
input GIN_257_171_gat;
input GIN_262_172_gat;
input GIN_263_173_gat;
input GIN_264_174_gat;
input GIN_265_175_gat;
input GIN_266_176_gat;
input GIN_267_177_gat;
input GIN_268_178_gat;
input GIN_269_179_gat;
input GIN_270_180_gat;
input GIN_271_181_gat;
input GIN_272_182_gat;
input GIN_273_183_gat;
input GIN_274_184_gat;
input GIN_275_185_gat;
input GIN_276_186_gat;
input GIN_277_187_gat;
input GIN_278_188_gat;
input GIN_279_189_gat;
input G452_190_gat;
input G483_191_gat;
input G543_192_gat;
input G559_193_gat;
input G567_194_gat;
input G651_195_gat;
input G661_196_gat;
input G860_197_gat;
input G868_198_gat;
input G1083_199_gat;
input G1341_200_gat;
input G1348_201_gat;
input G1384_202_gat;
input G1956_203_gat;
input G1961_204_gat;
input G1966_205_gat;
input G1971_206_gat;
input G1976_207_gat;
input G1981_208_gat;
input G1986_209_gat;
input G1991_210_gat;
input G1996_211_gat;
input G2066_212_gat;
input G2067_213_gat;
input G2072_214_gat;
input G2078_215_gat;
input G2084_216_gat;
input G2090_217_gat;
input G2096_218_gat;
input G2100_219_gat;
input G2104_220_gat;
input G2105_221_gat;
input G2106_222_gat;
input G2427_223_gat;
input G2430_224_gat;
input G2435_225_gat;
input G2438_226_gat;
input G2443_227_gat;
input G2446_228_gat;
input G2451_229_gat;
input G2454_230_gat;
input G2474_231_gat;
input G2678_232_gat;

output G169_114_gat;
output G174_115_gat;
output G177_116_gat;
output G178_117_gat;
output G179_118_gat;
output G180_119_gat;
output G181_120_gat;
output G182_121_gat;
output G183_122_gat;
output G184_123_gat;
output G185_124_gat;
output G186_125_gat;
output G189_126_gat;
output G190_127_gat;
output G191_128_gat;
output G192_129_gat;
output G193_130_gat;
output G194_131_gat;
output G195_132_gat;
output G196_133_gat;
output G197_134_gat;
output G198_135_gat;
output G199_136_gat;
output G200_137_gat;
output G201_138_gat;
output G202_139_gat;
output G203_140_gat;
output G204_141_gat;
output G205_142_gat;
output G206_143_gat;
output G207_144_gat;
output G208_145_gat;
output G209_146_gat;
output G210_147_gat;
output G211_148_gat;
output G212_149_gat;
output G213_150_gat;
output G214_151_gat;
output G215_152_gat;
output G239_153_gat;
output G240_154_gat;
output G241_155_gat;
output G242_156_gat;
output G243_157_gat;
output G244_158_gat;
output G245_159_gat;
output G246_160_gat;
output G247_161_gat;
output G248_162_gat;
output G249_163_gat;
output G250_164_gat;
output G251_165_gat;
output G252_166_gat;
output G253_167_gat;
output G254_168_gat;
output G255_169_gat;
output G256_170_gat;
output G257_171_gat;
output G262_172_gat;
output G263_173_gat;
output G264_174_gat;
output G265_175_gat;
output G266_176_gat;
output G267_177_gat;
output G268_178_gat;
output G269_179_gat;
output G270_180_gat;
output G271_181_gat;
output G272_182_gat;
output G273_183_gat;
output G274_184_gat;
output G275_185_gat;
output G276_186_gat;
output G277_187_gat;
output G278_188_gat;
output G279_189_gat;
output G350_301_gat;
output G335_299_gat;
output G409_298_gat;
output G369_289_gat;
output G367_288_gat;
output G411_264_gat;
output G337_263_gat;
output G384_262_gat;
output G218_311_gat;
output G219_302_gat;
output G220_306_gat;
output G221_305_gat;
output G235_307_gat;
output G236_303_gat;
output G237_309_gat;
output G238_304_gat;
output G158_349_gat;
output G259_414_gat;
output G391_379_gat;
output G173_389_gat;
output G223_413_gat;
output G234_376_gat;
output G217_423_gat;
output G325_507_gat;
output G261_506_gat;
output G319_656_gat;
output G160_609_gat;
output G162_612_gat;
output G164_607_gat;
output G166_625_gat;
output G168_623_gat;
output G171_621_gat;
output G153_671_gat;
output G176_803_gat;
output G188_761_gat;
output G299_692_gat;
output G301_694_gat;
output G286_696_gat;
output G303_698_gat;
output G288_700_gat;
output G305_702_gat;
output G290_704_gat;
output G284_847_gat;
output G321_848_gat;
output G297_849_gat;
output G280_850_gat;
output G148_851_gat;
output G282_922_gat;
output G323_923_gat;
output G156_1046_gat;
output G401_1276_gat;
output G227_1179_gat;
output G229_1180_gat;
output G311_1278_gat;
output G150_1277_gat;
output G145_1358_gat;
output G395_1392_gat;
output G295_1400_gat;
output G331_1401_gat;
output G397_1406_gat;
output G329_1414_gat;
output G231_1422_gat;
output G308_1425_gat;
output G225_1424_gat;

INVXL U_g1 (.A(G44_31_gat), .Y(G218_311_gat) );
INVXL U_g2 (.A(G132_105_gat), .Y(G219_302_gat) );
INVXL U_g3 (.A(G82_63_gat), .Y(G220_306_gat) );
INVXL U_g4 (.A(G96_75_gat), .Y(G221_305_gat) );
INVXL U_g5 (.A(G69_52_gat), .Y(G235_307_gat) );
INVXL U_g6 (.A(G120_95_gat), .Y(G236_303_gat) );
INVXL U_g7 (.A(G57_42_gat), .Y(G237_309_gat) );
INVXL U_g8 (.A(G108_85_gat), .Y(G238_304_gat) );
INVXL U_g9 (.A(G157_259_gat), .Y(G158_349_gat) );
INVXL U_g10 (.A(G258_321_gat), .Y(G259_414_gat) );
AND2XL U_g11 (.A(G391_379_gat), .B(G94_73_gat), .Y(G173_389_gat) );
INVXL U_g12 (.A(G1955_320_gat), .Y(G223_413_gat) );
OR2XL U_g13 (.A(G1955_320_ngat), .B(G567_194_ngat), .Y(G234_376_gat) );
INVXL U_g14 (.A(G216_333_gat), .Y(G217_423_gat) );
INVXL U_g15 (.A(G325_507_gat), .Y(G261_506_gat) );
INVXL U_g16 (.A(G1464_560_gat), .Y(G160_609_gat) );
INVXL U_g17 (.A(G1467_561_gat), .Y(G162_612_gat) );
INVXL U_g18 (.A(G1461_559_gat), .Y(G164_607_gat) );
INVXL U_g19 (.A(G1329_569_gat), .Y(G166_625_gat) );
INVXL U_g20 (.A(G1327_568_gat), .Y(G168_623_gat) );
INVXL U_g21 (.A(G857_567_gat), .Y(G171_621_gat) );
OR2XL U_g22 (.A(G152_599_gat), .B(G865_291_gat), .Y(G153_671_gat) );
INVXL U_g23 (.A(G175_710_gat), .Y(G176_803_gat) );
INVXL U_g24 (.A(G187_673_gat), .Y(G188_761_gat) );
OR2XL U_g25 (.A(G147_600_gat), .B(G146_758_gat), .Y(G148_851_gat) );
OR2XL U_g26 (.A(G155_967_ngat), .B(G154_964_ngat), .Y(G156_1046_gat) );
INVXL U_g27 (.A(G1830_1108_gat), .Y(G227_1179_gat) );
INVXL U_g28 (.A(G1553_1110_gat), .Y(G229_1180_gat) );
INVXL U_g29 (.A(G311_1278_gat), .Y(G150_1277_gat) );
OR2XL U_g30 (.A(G144_601_gat), .B(G143_1330_gat), .Y(G145_1358_gat) );
INVXL U_g31 (.A(G473_1420_gat), .Y(G231_1422_gat) );
INVXL U_g32 (.A(G308_1425_gat), .Y(G225_1424_gat) );
INVXL U_g33 (.A(G2678_232_gat), .Y(G2682_233_gat) );
INVXL U_g34 (.A(G2474_231_gat), .Y(G2478_234_gat) );
INVXL U_g35 (.A(G2454_230_gat), .Y(G2458_235_gat) );
INVXL U_g36 (.A(G2451_229_gat), .Y(G2457_236_gat) );
INVXL U_g37 (.A(G2446_228_gat), .Y(G2450_237_gat) );
INVXL U_g38 (.A(G2443_227_gat), .Y(G2449_238_gat) );
INVXL U_g39 (.A(G2438_226_gat), .Y(G2442_239_gat) );
INVXL U_g40 (.A(G2435_225_gat), .Y(G2441_240_gat) );
INVXL U_g41 (.A(G2430_224_gat), .Y(G2434_241_gat) );
INVXL U_g42 (.A(G2427_223_gat), .Y(G2433_242_gat) );
BUFX20 U_g43 (.A(G2105_221_gat), .Y(G1655_243_gat) );
BUFX20 U_g44 (.A(G2105_221_gat), .Y(G1418_244_gat) );
BUFX20 U_g45 (.A(G2104_220_gat), .Y(G1631_245_gat) );
BUFX20 U_g46 (.A(G2104_220_gat), .Y(G1394_246_gat) );
INVXL U_g47 (.A(G2100_219_gat), .Y(G2103_247_gat) );
BUFX20 U_g48 (.A(G2100_219_gat), .Y(G2699_248_gat) );
INVXL U_g49 (.A(G2096_218_gat), .Y(G2099_249_gat) );
BUFX20 U_g50 (.A(G2096_218_gat), .Y(G2702_250_gat) );
INVXL U_g51 (.A(G2090_217_gat), .Y(G2094_251_gat) );
BUFX20 U_g52 (.A(G2090_217_gat), .Y(G2691_252_gat) );
INVXL U_g53 (.A(G2084_216_gat), .Y(G2088_253_gat) );
BUFX20 U_g54 (.A(G2084_216_gat), .Y(G2694_254_gat) );
INVXL U_g55 (.A(G2078_215_gat), .Y(G2082_255_gat) );
BUFX20 U_g56 (.A(G2078_215_gat), .Y(G2683_256_gat) );
INVXL U_g57 (.A(G2072_214_gat), .Y(G2076_257_gat) );
BUFX20 U_g58 (.A(G2072_214_gat), .Y(G2686_258_gat) );
AND4XL U_g59 (.A(G2072_214_gat), .B(G2078_215_gat), .C(G2084_216_gat), .D(G2090_217_gat), .Y(G157_259_gat) );
INVXL U_g60 (.A(G2067_213_gat), .Y(G2070_260_gat) );
BUFX20 U_g61 (.A(G2067_213_gat), .Y(G2675_261_gat) );
INVXL U_g62 (.A(G1996_211_gat), .Y(G1999_265_gat) );
BUFX20 U_g63 (.A(G1996_211_gat), .Y(G2505_266_gat) );
INVXL U_g64 (.A(G1991_210_gat), .Y(G1994_267_gat) );
BUFX20 U_g65 (.A(G1991_210_gat), .Y(G2508_268_gat) );
INVXL U_g66 (.A(G1986_209_gat), .Y(G1989_269_gat) );
BUFX20 U_g67 (.A(G1986_209_gat), .Y(G2495_270_gat) );
INVXL U_g68 (.A(G1981_208_gat), .Y(G1984_271_gat) );
BUFX20 U_g69 (.A(G1981_208_gat), .Y(G2498_272_gat) );
INVXL U_g70 (.A(G1976_207_gat), .Y(G1979_273_gat) );
BUFX20 U_g71 (.A(G1976_207_gat), .Y(G2487_274_gat) );
INVXL U_g72 (.A(G1971_206_gat), .Y(G1974_275_gat) );
BUFX20 U_g73 (.A(G1971_206_gat), .Y(G2490_276_gat) );
INVXL U_g74 (.A(G1966_205_gat), .Y(G1969_277_gat) );
BUFX20 U_g75 (.A(G1966_205_gat), .Y(G2479_278_gat) );
INVXL U_g76 (.A(G1961_204_gat), .Y(G1964_279_gat) );
BUFX20 U_g77 (.A(G1961_204_gat), .Y(G2482_280_gat) );
INVXL U_g78 (.A(G1956_203_gat), .Y(G1959_281_gat) );
BUFX20 U_g79 (.A(G1956_203_gat), .Y(G2471_282_gat) );
INVXL U_g80 (.A(G1384_202_gat), .Y(G1385_283_gat) );
INVXL U_g81 (.A(G1348_201_gat), .Y(G1351_284_gat) );
BUFX20 U_g82 (.A(G1348_201_gat), .Y(G2461_285_gat) );
INVXL U_g83 (.A(G1341_200_gat), .Y(G1344_286_gat) );
BUFX20 U_g84 (.A(G1341_200_gat), .Y(G2464_287_gat) );
INVXL U_g85 (.A(G868_198_gat), .Y(G875_290_gat) );
INVXL U_g86 (.A(G860_197_gat), .Y(G865_291_gat) );
BUFX20 U_g87 (.A(G661_196_gat), .Y(G480_292_gat) );
BUFX20 U_g88 (.A(G651_195_gat), .Y(G1284_293_gat) );
BUFX20 U_g89 (.A(G651_195_gat), .Y(G795_294_gat) );
INVXL U_g90 (.A(G559_193_gat), .Y(G560_295_gat) );
BUFX20 U_g91 (.A(G543_192_gat), .Y(G1261_296_gat) );
BUFX20 U_g92 (.A(G543_192_gat), .Y(G772_297_gat) );
BUFX20 U_g93 (.A(G452_190_gat), .Y(G391_379_gat) );
AND4XL U_g94 (.A(G69_52_gat), .B(G108_85_gat), .C(G57_42_gat), .D(G120_95_gat), .Y(G1254_308_gat) );
AND4XL U_g95 (.A(G44_31_gat), .B(G96_75_gat), .C(G82_63_gat), .D(G132_105_gat), .Y(G1251_310_gat) );
BUFX20 U_g96 (.A(G37_28_gat), .Y(G486_312_gat) );
BUFX20 U_g97 (.A(G29_22_gat), .Y(G2012_313_gat) );
BUFX20 U_g98 (.A(G29_22_gat), .Y(G2001_314_gat) );
BUFX20 U_g99 (.A(G16_11_gat), .Y(G1721_315_gat) );
BUFX20 U_g100 (.A(G16_11_gat), .Y(G1710_316_gat) );
AND2XL U_g101 (.A(G868_198_gat), .B(G11_8_gat), .Y(G882_317_gat) );
BUFX20 U_g102 (.A(G8_7_gat), .Y(G658_318_gat) );
BUFX20 U_g103 (.A(G8_7_gat), .Y(G655_319_gat) );
AND2XL U_g104 (.A(G661_196_gat), .B(G7_6_gat), .Y(G1955_320_gat) );
AND3XL U_g105 (.A(G661_196_gat), .B(G15_10_gat), .C(G2_1_gat), .Y(G258_321_gat) );
AND2XL U_g106 (.A(G3_2_gat), .B(G1_0_gat), .Y(G546_322_gat) );
OR2XL U_g107 (.A(G2682_233_ngat), .B(G2675_261_ngat), .Y(G1776_323_gat) );
OR2XL U_g108 (.A(G2478_234_ngat), .B(G2471_282_ngat), .Y(G1499_324_gat) );
OR2XL U_g109 (.A(G2457_236_ngat), .B(G2454_230_ngat), .Y(G2459_325_gat) );
OR2XL U_g110 (.A(G2458_235_ngat), .B(G2451_229_ngat), .Y(G2460_326_gat) );
OR2XL U_g111 (.A(G2449_238_ngat), .B(G2446_228_ngat), .Y(G1493_327_gat) );
OR2XL U_g112 (.A(G2450_237_ngat), .B(G2443_227_ngat), .Y(G1494_328_gat) );
OR2XL U_g113 (.A(G2441_240_ngat), .B(G2438_226_ngat), .Y(G1484_329_gat) );
OR2XL U_g114 (.A(G2442_239_ngat), .B(G2435_225_ngat), .Y(G1485_330_gat) );
OR2XL U_g115 (.A(G2433_242_ngat), .B(G2430_224_ngat), .Y(G1475_331_gat) );
OR2XL U_g116 (.A(G2434_241_ngat), .B(G2427_223_ngat), .Y(G1476_332_gat) );
AND2XL U_g117 (.A(G1955_320_gat), .B(G2106_222_gat), .Y(G216_333_gat) );
INVXL U_g118 (.A(G1655_243_gat), .Y(G1667_334_gat) );
AND2XL U_g119 (.A(G1418_244_gat), .B(G1394_246_gat), .Y(G1460_335_gat) );
INVXL U_g120 (.A(G1418_244_gat), .Y(G1430_336_gat) );
INVXL U_g121 (.A(G1631_245_gat), .Y(G1643_337_gat) );
INVXL U_g122 (.A(G1394_246_gat), .Y(G1406_338_gat) );
INVXL U_g123 (.A(G2699_248_gat), .Y(G2705_339_gat) );
INVXL U_g124 (.A(G2702_250_gat), .Y(G2706_340_gat) );
BUFX20 U_g125 (.A(G2094_251_gat), .Y(G2775_341_gat) );
INVXL U_g126 (.A(G2691_252_gat), .Y(G2697_342_gat) );
BUFX20 U_g127 (.A(G2088_253_gat), .Y(G2767_343_gat) );
INVXL U_g128 (.A(G2694_254_gat), .Y(G2698_344_gat) );
BUFX20 U_g129 (.A(G2082_255_gat), .Y(G2759_345_gat) );
INVXL U_g130 (.A(G2683_256_gat), .Y(G2689_346_gat) );
BUFX20 U_g131 (.A(G2076_257_gat), .Y(G2751_347_gat) );
INVXL U_g132 (.A(G2686_258_gat), .Y(G2690_348_gat) );
BUFX20 U_g133 (.A(G2070_260_gat), .Y(G2743_350_gat) );
INVXL U_g134 (.A(G2675_261_gat), .Y(G2681_351_gat) );
BUFX20 U_g135 (.A(G1999_265_gat), .Y(G2735_352_gat) );
INVXL U_g136 (.A(G2505_266_gat), .Y(G2511_353_gat) );
BUFX20 U_g137 (.A(G1994_267_gat), .Y(G2623_354_gat) );
INVXL U_g138 (.A(G2508_268_gat), .Y(G2512_355_gat) );
BUFX20 U_g139 (.A(G1989_269_gat), .Y(G2615_356_gat) );
INVXL U_g140 (.A(G2495_270_gat), .Y(G2501_357_gat) );
BUFX20 U_g141 (.A(G1984_271_gat), .Y(G2607_358_gat) );
INVXL U_g142 (.A(G2498_272_gat), .Y(G2502_359_gat) );
BUFX20 U_g143 (.A(G1979_273_gat), .Y(G2599_360_gat) );
INVXL U_g144 (.A(G2487_274_gat), .Y(G2493_361_gat) );
BUFX20 U_g145 (.A(G1974_275_gat), .Y(G2591_362_gat) );
INVXL U_g146 (.A(G2490_276_gat), .Y(G2494_363_gat) );
BUFX20 U_g147 (.A(G1969_277_gat), .Y(G2583_364_gat) );
INVXL U_g148 (.A(G2479_278_gat), .Y(G2485_365_gat) );
BUFX20 U_g149 (.A(G1964_279_gat), .Y(G2575_366_gat) );
INVXL U_g150 (.A(G2482_280_gat), .Y(G2486_367_gat) );
BUFX20 U_g151 (.A(G1959_281_gat), .Y(G2567_368_gat) );
INVXL U_g152 (.A(G2471_282_gat), .Y(G2477_369_gat) );
BUFX20 U_g153 (.A(G1351_284_gat), .Y(G2559_370_gat) );
INVXL U_g154 (.A(G2461_285_gat), .Y(G2467_371_gat) );
BUFX20 U_g155 (.A(G1344_286_gat), .Y(G2551_372_gat) );
INVXL U_g156 (.A(G2464_287_gat), .Y(G2468_373_gat) );
INVXL U_g157 (.A(G1284_293_gat), .Y(G1296_374_gat) );
INVXL U_g158 (.A(G795_294_gat), .Y(G807_375_gat) );
INVXL U_g159 (.A(G1261_296_gat), .Y(G1273_377_gat) );
INVXL U_g160 (.A(G772_297_gat), .Y(G784_378_gat) );
AND3XL U_g161 (.A(G1655_243_gat), .B(G1631_245_gat), .C(G118_93_gat), .Y(G1681_380_gat) );
AND3XL U_g162 (.A(G1655_243_gat), .B(G1631_245_gat), .C(G117_92_gat), .Y(G1689_381_gat) );
AND3XL U_g163 (.A(G1655_243_gat), .B(G1631_245_gat), .C(G116_91_gat), .Y(G1693_382_gat) );
AND3XL U_g164 (.A(G1655_243_gat), .B(G1631_245_gat), .C(G115_90_gat), .Y(G1697_383_gat) );
AND3XL U_g165 (.A(G1418_244_gat), .B(G1394_246_gat), .C(G114_89_gat), .Y(G1444_384_gat) );
AND3XL U_g166 (.A(G1418_244_gat), .B(G1394_246_gat), .C(G113_88_gat), .Y(G1448_385_gat) );
AND3XL U_g167 (.A(G1418_244_gat), .B(G1394_246_gat), .C(G112_87_gat), .Y(G1452_386_gat) );
AND3XL U_g168 (.A(G1418_244_gat), .B(G1394_246_gat), .C(G111_86_gat), .Y(G1456_387_gat) );
AND3XL U_g169 (.A(G1655_243_gat), .B(G1631_245_gat), .C(G107_84_gat), .Y(G1685_388_gat) );
AND3XL U_g170 (.A(G795_294_gat), .B(G772_297_gat), .C(G80_61_gat), .Y(G821_390_gat) );
AND3XL U_g171 (.A(G795_294_gat), .B(G772_297_gat), .C(G79_60_gat), .Y(G829_391_gat) );
AND3XL U_g172 (.A(G795_294_gat), .B(G772_297_gat), .C(G78_59_gat), .Y(G833_392_gat) );
AND3XL U_g173 (.A(G795_294_gat), .B(G772_297_gat), .C(G77_58_gat), .Y(G837_393_gat) );
AND3XL U_g174 (.A(G1284_293_gat), .B(G1261_296_gat), .C(G76_57_gat), .Y(G1310_394_gat) );
AND3XL U_g175 (.A(G1284_293_gat), .B(G1261_296_gat), .C(G75_56_gat), .Y(G1314_395_gat) );
AND3XL U_g176 (.A(G1284_293_gat), .B(G1261_296_gat), .C(G74_55_gat), .Y(G1318_396_gat) );
AND3XL U_g177 (.A(G1284_293_gat), .B(G1261_296_gat), .C(G73_54_gat), .Y(G1322_397_gat) );
AND3XL U_g178 (.A(G1284_293_gat), .B(G1261_296_gat), .C(G72_53_gat), .Y(G1326_398_gat) );
AND3XL U_g179 (.A(G795_294_gat), .B(G772_297_gat), .C(G68_51_gat), .Y(G825_399_gat) );
AND2XL U_g180 (.A(G1251_310_gat), .B(G1254_308_gat), .Y(G325_507_gat) );
INVXL U_g181 (.A(G1254_308_gat), .Y(G1256_401_gat) );
INVXL U_g182 (.A(G1251_310_gat), .Y(G1253_402_gat) );
INVXL U_g183 (.A(G486_312_gat), .Y(G487_403_gat) );
INVXL U_g184 (.A(G2012_313_gat), .Y(G2018_404_gat) );
INVXL U_g185 (.A(G2001_314_gat), .Y(G2007_405_gat) );
INVXL U_g186 (.A(G1721_315_gat), .Y(G1728_406_gat) );
INVXL U_g187 (.A(G1710_316_gat), .Y(G1716_407_gat) );
AND2XL U_g188 (.A(G875_290_gat), .B(G11_8_gat), .Y(G881_408_gat) );
BUFX20 U_g189 (.A(G658_318_gat), .Y(G1831_409_gat) );
BUFX20 U_g190 (.A(G658_318_gat), .Y(G1893_410_gat) );
BUFX20 U_g191 (.A(G655_319_gat), .Y(G748_411_gat) );
BUFX20 U_g192 (.A(G655_319_gat), .Y(G994_412_gat) );
INVXL U_g193 (.A(G546_322_gat), .Y(G547_415_gat) );
OR2XL U_g194 (.A(G2681_351_ngat), .B(G2678_232_ngat), .Y(G1775_416_gat) );
OR2XL U_g195 (.A(G2477_369_ngat), .B(G2474_231_ngat), .Y(G1498_417_gat) );
OR2XL U_g196 (.A(G2460_326_ngat), .B(G2459_325_ngat), .Y(G2518_418_gat) );
OR2XL U_g197 (.A(G1494_328_ngat), .B(G1493_327_ngat), .Y(G1495_419_gat) );
OR2XL U_g198 (.A(G1485_330_ngat), .B(G1484_329_ngat), .Y(G1486_420_gat) );
OR2XL U_g199 (.A(G1476_332_ngat), .B(G1475_331_ngat), .Y(G1477_421_gat) );
AND2XL U_g200 (.A(G1253_402_gat), .B(G2106_222_gat), .Y(G550_422_gat) );
AND2XL U_g201 (.A(G1418_244_gat), .B(G1406_338_gat), .Y(G1459_424_gat) );
AND2XL U_g202 (.A(G1430_336_gat), .B(G1406_338_gat), .Y(G1457_425_gat) );
AND2XL U_g203 (.A(G1430_336_gat), .B(G1394_246_gat), .Y(G1458_426_gat) );
OR2XL U_g204 (.A(G2706_340_ngat), .B(G2699_248_ngat), .Y(G2708_427_gat) );
OR2XL U_g205 (.A(G2705_339_ngat), .B(G2702_250_ngat), .Y(G2707_428_gat) );
INVXL U_g206 (.A(G2775_341_gat), .Y(G2781_429_gat) );
OR2XL U_g207 (.A(G2698_344_ngat), .B(G2691_252_ngat), .Y(G1794_430_gat) );
INVXL U_g208 (.A(G2767_343_gat), .Y(G2773_431_gat) );
OR2XL U_g209 (.A(G2697_342_ngat), .B(G2694_254_ngat), .Y(G1793_432_gat) );
INVXL U_g210 (.A(G2759_345_gat), .Y(G2765_433_gat) );
OR2XL U_g211 (.A(G2690_348_ngat), .B(G2683_256_ngat), .Y(G1785_434_gat) );
INVXL U_g212 (.A(G2751_347_gat), .Y(G2757_435_gat) );
OR2XL U_g213 (.A(G2689_346_ngat), .B(G2686_258_ngat), .Y(G1784_436_gat) );
INVXL U_g214 (.A(G2743_350_gat), .Y(G2749_437_gat) );
INVXL U_g215 (.A(G2735_352_gat), .Y(G2741_438_gat) );
OR2XL U_g216 (.A(G2512_355_ngat), .B(G2505_266_ngat), .Y(G2514_439_gat) );
INVXL U_g217 (.A(G2623_354_gat), .Y(G2629_440_gat) );
OR2XL U_g218 (.A(G2511_353_ngat), .B(G2508_268_ngat), .Y(G2513_441_gat) );
INVXL U_g219 (.A(G2615_356_gat), .Y(G2621_442_gat) );
OR2XL U_g220 (.A(G2502_359_ngat), .B(G2495_270_ngat), .Y(G2504_443_gat) );
INVXL U_g221 (.A(G2607_358_gat), .Y(G2613_444_gat) );
OR2XL U_g222 (.A(G2501_357_ngat), .B(G2498_272_ngat), .Y(G2503_445_gat) );
INVXL U_g223 (.A(G2599_360_gat), .Y(G2605_446_gat) );
OR2XL U_g224 (.A(G2494_363_ngat), .B(G2487_274_ngat), .Y(G1517_447_gat) );
INVXL U_g225 (.A(G2591_362_gat), .Y(G2597_448_gat) );
OR2XL U_g226 (.A(G2493_361_ngat), .B(G2490_276_ngat), .Y(G1516_449_gat) );
INVXL U_g227 (.A(G2583_364_gat), .Y(G2589_450_gat) );
OR2XL U_g228 (.A(G2486_367_ngat), .B(G2479_278_ngat), .Y(G1508_451_gat) );
INVXL U_g229 (.A(G2575_366_gat), .Y(G2581_452_gat) );
OR2XL U_g230 (.A(G2485_365_ngat), .B(G2482_280_ngat), .Y(G1507_453_gat) );
INVXL U_g231 (.A(G2567_368_gat), .Y(G2573_454_gat) );
INVXL U_g232 (.A(G2559_370_gat), .Y(G2565_455_gat) );
OR2XL U_g233 (.A(G2468_373_ngat), .B(G2461_285_ngat), .Y(G2470_456_gat) );
INVXL U_g234 (.A(G2551_372_gat), .Y(G2557_457_gat) );
OR2XL U_g235 (.A(G2467_371_ngat), .B(G2464_287_ngat), .Y(G2469_458_gat) );
AND2XL U_g236 (.A(G1284_293_gat), .B(G1273_377_gat), .Y(G1317_459_gat) );
AND2XL U_g237 (.A(G1256_401_gat), .B(G567_194_gat), .Y(G552_460_gat) );
AND3XL U_g238 (.A(G1667_334_gat), .B(G1643_337_gat), .C(G142_113_gat), .Y(G1678_461_gat) );
AND3XL U_g239 (.A(G1667_334_gat), .B(G1643_337_gat), .C(G141_112_gat), .Y(G1686_462_gat) );
AND3XL U_g240 (.A(G1667_334_gat), .B(G1643_337_gat), .C(G140_111_gat), .Y(G1690_463_gat) );
AND3XL U_g241 (.A(G1667_334_gat), .B(G1643_337_gat), .C(G139_110_gat), .Y(G1694_464_gat) );
AND3XL U_g242 (.A(G1430_336_gat), .B(G1406_338_gat), .C(G138_109_gat), .Y(G1441_465_gat) );
AND3XL U_g243 (.A(G1430_336_gat), .B(G1406_338_gat), .C(G137_108_gat), .Y(G1445_466_gat) );
AND3XL U_g244 (.A(G1430_336_gat), .B(G1406_338_gat), .C(G136_107_gat), .Y(G1449_467_gat) );
AND3XL U_g245 (.A(G1430_336_gat), .B(G1406_338_gat), .C(G135_106_gat), .Y(G1453_468_gat) );
AND3XL U_g246 (.A(G1667_334_gat), .B(G1643_337_gat), .C(G131_104_gat), .Y(G1682_469_gat) );
AND3XL U_g247 (.A(G1655_243_gat), .B(G1643_337_gat), .C(G130_103_gat), .Y(G1680_470_gat) );
AND3XL U_g248 (.A(G1655_243_gat), .B(G1643_337_gat), .C(G129_102_gat), .Y(G1688_471_gat) );
AND3XL U_g249 (.A(G1655_243_gat), .B(G1643_337_gat), .C(G128_101_gat), .Y(G1692_472_gat) );
AND3XL U_g250 (.A(G1655_243_gat), .B(G1643_337_gat), .C(G127_100_gat), .Y(G1696_473_gat) );
AND3XL U_g251 (.A(G1418_244_gat), .B(G1406_338_gat), .C(G126_99_gat), .Y(G1443_474_gat) );
AND3XL U_g252 (.A(G1418_244_gat), .B(G1406_338_gat), .C(G125_98_gat), .Y(G1447_475_gat) );
AND3XL U_g253 (.A(G1418_244_gat), .B(G1406_338_gat), .C(G124_97_gat), .Y(G1451_476_gat) );
AND3XL U_g254 (.A(G1418_244_gat), .B(G1406_338_gat), .C(G123_96_gat), .Y(G1455_477_gat) );
AND3XL U_g255 (.A(G1655_243_gat), .B(G1643_337_gat), .C(G119_94_gat), .Y(G1684_478_gat) );
AND3XL U_g256 (.A(G1667_334_gat), .B(G1631_245_gat), .C(G106_83_gat), .Y(G1679_479_gat) );
AND3XL U_g257 (.A(G1667_334_gat), .B(G1631_245_gat), .C(G105_82_gat), .Y(G1687_480_gat) );
AND3XL U_g258 (.A(G1667_334_gat), .B(G1631_245_gat), .C(G104_81_gat), .Y(G1691_481_gat) );
AND3XL U_g259 (.A(G1667_334_gat), .B(G1631_245_gat), .C(G103_80_gat), .Y(G1695_482_gat) );
AND3XL U_g260 (.A(G1430_336_gat), .B(G1394_246_gat), .C(G102_79_gat), .Y(G1442_483_gat) );
AND3XL U_g261 (.A(G1430_336_gat), .B(G1394_246_gat), .C(G101_78_gat), .Y(G1446_484_gat) );
AND3XL U_g262 (.A(G1430_336_gat), .B(G1394_246_gat), .C(G100_77_gat), .Y(G1450_485_gat) );
AND3XL U_g263 (.A(G1430_336_gat), .B(G1394_246_gat), .C(G99_76_gat), .Y(G1454_486_gat) );
AND3XL U_g264 (.A(G1667_334_gat), .B(G1631_245_gat), .C(G95_74_gat), .Y(G1683_487_gat) );
AND3XL U_g265 (.A(G807_375_gat), .B(G784_378_gat), .C(G93_72_gat), .Y(G818_488_gat) );
AND3XL U_g266 (.A(G807_375_gat), .B(G784_378_gat), .C(G92_71_gat), .Y(G826_489_gat) );
AND3XL U_g267 (.A(G807_375_gat), .B(G784_378_gat), .C(G91_70_gat), .Y(G830_490_gat) );
AND3XL U_g268 (.A(G807_375_gat), .B(G784_378_gat), .C(G90_69_gat), .Y(G834_491_gat) );
AND3XL U_g269 (.A(G1296_374_gat), .B(G1273_377_gat), .C(G89_68_gat), .Y(G1307_492_gat) );
AND3XL U_g270 (.A(G1296_374_gat), .B(G1273_377_gat), .C(G88_67_gat), .Y(G1311_493_gat) );
AND3XL U_g271 (.A(G1296_374_gat), .B(G1273_377_gat), .C(G87_66_gat), .Y(G1315_494_gat) );
AND3XL U_g272 (.A(G1296_374_gat), .B(G1273_377_gat), .C(G86_65_gat), .Y(G1319_495_gat) );
AND3XL U_g273 (.A(G1296_374_gat), .B(G1273_377_gat), .C(G85_64_gat), .Y(G1323_496_gat) );
AND3XL U_g274 (.A(G807_375_gat), .B(G784_378_gat), .C(G81_62_gat), .Y(G822_497_gat) );
AND3XL U_g275 (.A(G795_294_gat), .B(G784_378_gat), .C(G67_50_gat), .Y(G820_498_gat) );
AND3XL U_g276 (.A(G795_294_gat), .B(G784_378_gat), .C(G66_49_gat), .Y(G828_499_gat) );
AND3XL U_g277 (.A(G795_294_gat), .B(G784_378_gat), .C(G65_48_gat), .Y(G832_500_gat) );
AND3XL U_g278 (.A(G795_294_gat), .B(G784_378_gat), .C(G64_47_gat), .Y(G836_501_gat) );
AND3XL U_g279 (.A(G1284_293_gat), .B(G1273_377_gat), .C(G63_46_gat), .Y(G1309_502_gat) );
AND3XL U_g280 (.A(G1284_293_gat), .B(G1273_377_gat), .C(G62_45_gat), .Y(G1313_503_gat) );
AND3XL U_g281 (.A(G1284_293_gat), .B(G1273_377_gat), .C(G61_44_gat), .Y(G1321_504_gat) );
AND3XL U_g282 (.A(G1284_293_gat), .B(G1273_377_gat), .C(G60_43_gat), .Y(G1325_505_gat) );
AND3XL U_g283 (.A(G795_294_gat), .B(G784_378_gat), .C(G56_41_gat), .Y(G824_508_gat) );
AND3XL U_g284 (.A(G807_375_gat), .B(G772_297_gat), .C(G55_40_gat), .Y(G819_509_gat) );
AND3XL U_g285 (.A(G807_375_gat), .B(G772_297_gat), .C(G54_39_gat), .Y(G827_510_gat) );
AND3XL U_g286 (.A(G807_375_gat), .B(G772_297_gat), .C(G53_38_gat), .Y(G831_511_gat) );
AND3XL U_g287 (.A(G807_375_gat), .B(G772_297_gat), .C(G52_37_gat), .Y(G835_512_gat) );
AND3XL U_g288 (.A(G1296_374_gat), .B(G1261_296_gat), .C(G51_36_gat), .Y(G1308_513_gat) );
AND3XL U_g289 (.A(G1296_374_gat), .B(G1261_296_gat), .C(G50_35_gat), .Y(G1312_514_gat) );
AND3XL U_g290 (.A(G1296_374_gat), .B(G1261_296_gat), .C(G49_34_gat), .Y(G1316_515_gat) );
AND3XL U_g291 (.A(G1296_374_gat), .B(G1261_296_gat), .C(G48_33_gat), .Y(G1320_516_gat) );
AND3XL U_g292 (.A(G1296_374_gat), .B(G1261_296_gat), .C(G47_32_gat), .Y(G1324_517_gat) );
AND3XL U_g293 (.A(G807_375_gat), .B(G772_297_gat), .C(G43_30_gat), .Y(G823_518_gat) );
AND2XL U_g294 (.A(G2018_404_gat), .B(G35_26_gat), .Y(G2035_519_gat) );
AND2XL U_g295 (.A(G2018_404_gat), .B(G34_25_gat), .Y(G2033_520_gat) );
AND2XL U_g296 (.A(G2007_405_gat), .B(G33_24_gat), .Y(G2029_521_gat) );
AND2XL U_g297 (.A(G2007_405_gat), .B(G32_23_gat), .Y(G2025_522_gat) );
AND2XL U_g298 (.A(G2018_404_gat), .B(G28_21_gat), .Y(G2037_523_gat) );
AND2XL U_g299 (.A(G2018_404_gat), .B(G27_20_gat), .Y(G2031_524_gat) );
AND2XL U_g300 (.A(G2007_405_gat), .B(G26_19_gat), .Y(G2027_525_gat) );
AND2XL U_g301 (.A(G2007_405_gat), .B(G25_18_gat), .Y(G2023_526_gat) );
AND2XL U_g302 (.A(G1728_406_gat), .B(G24_17_gat), .Y(G1750_527_gat) );
AND2XL U_g303 (.A(G1728_406_gat), .B(G23_16_gat), .Y(G1746_528_gat) );
AND2XL U_g304 (.A(G1728_406_gat), .B(G22_15_gat), .Y(G1744_529_gat) );
AND2XL U_g305 (.A(G1728_406_gat), .B(G21_14_gat), .Y(G1742_530_gat) );
AND2XL U_g306 (.A(G1716_407_gat), .B(G20_13_gat), .Y(G1738_531_gat) );
AND2XL U_g307 (.A(G1716_407_gat), .B(G19_12_gat), .Y(G1734_532_gat) );
OR2XL U_g308 (.A(G882_317_gat), .B(G881_408_gat), .Y(G894_533_gat) );
AND2XL U_g309 (.A(G1728_406_gat), .B(G6_5_gat), .Y(G1748_534_gat) );
AND2XL U_g310 (.A(G1716_407_gat), .B(G5_4_gat), .Y(G1740_535_gat) );
AND2XL U_g311 (.A(G1716_407_gat), .B(G4_3_gat), .Y(G1736_536_gat) );
OR2XL U_g312 (.A(G1776_323_ngat), .B(G1775_416_ngat), .Y(G1777_537_gat) );
OR2XL U_g313 (.A(G1499_324_ngat), .B(G1498_417_ngat), .Y(G1500_538_gat) );
INVXL U_g314 (.A(G2518_418_gat), .Y(G2522_539_gat) );
BUFX20 U_g315 (.A(G1495_419_gat), .Y(G1525_540_gat) );
BUFX20 U_g316 (.A(G1495_419_gat), .Y(G1521_541_gat) );
INVXL U_g317 (.A(G1486_420_gat), .Y(G1490_542_gat) );
INVXL U_g318 (.A(G1477_421_gat), .Y(G1481_543_gat) );
INVXL U_g319 (.A(G550_422_gat), .Y(G551_544_gat) );
OR4XL U_g320 (.A(G1460_335_gat), .B(G1459_424_gat), .C(G1458_426_gat), .D(G1457_425_gat), .Y(G1473_545_gat) );
OR2XL U_g321 (.A(G2708_427_ngat), .B(G2707_428_ngat), .Y(G2730_546_gat) );
OR2XL U_g322 (.A(G1794_430_ngat), .B(G1793_432_ngat), .Y(G1795_547_gat) );
OR2XL U_g323 (.A(G1785_434_ngat), .B(G1784_436_ngat), .Y(G1786_548_gat) );
OR2XL U_g324 (.A(G2514_439_ngat), .B(G2513_441_ngat), .Y(G2525_549_gat) );
OR2XL U_g325 (.A(G2504_443_ngat), .B(G2503_445_ngat), .Y(G2528_550_gat) );
OR2XL U_g326 (.A(G1517_447_ngat), .B(G1516_449_ngat), .Y(G1518_551_gat) );
OR2XL U_g327 (.A(G1508_451_ngat), .B(G1507_453_ngat), .Y(G1509_552_gat) );
OR2XL U_g328 (.A(G2470_456_ngat), .B(G2469_458_ngat), .Y(G2515_553_gat) );
INVXL U_g329 (.A(G552_460_gat), .Y(G553_554_gat) );
OR4XL U_g330 (.A(G1681_380_gat), .B(G1680_470_gat), .C(G1679_479_gat), .D(G1678_461_gat), .Y(G2634_555_gat) );
OR4XL U_g331 (.A(G1689_381_gat), .B(G1688_471_gat), .C(G1687_480_gat), .D(G1686_462_gat), .Y(G1701_556_gat) );
OR4XL U_g332 (.A(G1693_382_gat), .B(G1692_472_gat), .C(G1691_481_gat), .D(G1690_463_gat), .Y(G1704_557_gat) );
OR4XL U_g333 (.A(G1697_383_gat), .B(G1696_473_gat), .C(G1695_482_gat), .D(G1694_464_gat), .Y(G1707_558_gat) );
OR4XL U_g334 (.A(G1444_384_gat), .B(G1443_474_gat), .C(G1442_483_gat), .D(G1441_465_gat), .Y(G1461_559_gat) );
OR4XL U_g335 (.A(G1448_385_gat), .B(G1447_475_gat), .C(G1446_484_gat), .D(G1445_466_gat), .Y(G1464_560_gat) );
OR4XL U_g336 (.A(G1452_386_gat), .B(G1451_476_gat), .C(G1450_485_gat), .D(G1449_467_gat), .Y(G1467_561_gat) );
OR4XL U_g337 (.A(G1456_387_gat), .B(G1455_477_gat), .C(G1454_486_gat), .D(G1453_468_gat), .Y(G1470_562_gat) );
OR4XL U_g338 (.A(G1685_388_gat), .B(G1684_478_gat), .C(G1683_487_gat), .D(G1682_469_gat), .Y(G1698_563_gat) );
OR4XL U_g339 (.A(G821_390_gat), .B(G820_498_gat), .C(G819_509_gat), .D(G818_488_gat), .Y(G838_564_gat) );
OR4XL U_g340 (.A(G829_391_gat), .B(G828_499_gat), .C(G827_510_gat), .D(G826_489_gat), .Y(G846_565_gat) );
OR4XL U_g341 (.A(G833_392_gat), .B(G832_500_gat), .C(G831_511_gat), .D(G830_490_gat), .Y(G854_566_gat) );
OR4XL U_g342 (.A(G837_393_gat), .B(G836_501_gat), .C(G835_512_gat), .D(G834_491_gat), .Y(G857_567_gat) );
OR4XL U_g343 (.A(G1310_394_gat), .B(G1309_502_gat), .C(G1308_513_gat), .D(G1307_492_gat), .Y(G1327_568_gat) );
OR4XL U_g344 (.A(G1314_395_gat), .B(G1313_503_gat), .C(G1312_514_gat), .D(G1311_493_gat), .Y(G1329_569_gat) );
OR4XL U_g345 (.A(G1318_396_gat), .B(G1317_459_gat), .C(G1316_515_gat), .D(G1315_494_gat), .Y(G1331_570_gat) );
OR4XL U_g346 (.A(G1322_397_gat), .B(G1321_504_gat), .C(G1320_516_gat), .D(G1319_495_gat), .Y(G1333_571_gat) );
OR4XL U_g347 (.A(G1326_398_gat), .B(G1325_505_gat), .C(G1324_517_gat), .D(G1323_496_gat), .Y(G1335_572_gat) );
OR4XL U_g348 (.A(G825_399_gat), .B(G824_508_gat), .C(G823_518_gat), .D(G822_497_gat), .Y(G841_573_gat) );
INVXL U_g349 (.A(G1777_537_gat), .Y(G1781_574_gat) );
INVXL U_g350 (.A(G1500_538_gat), .Y(G1504_575_gat) );
OR2XL U_g351 (.A(G2522_539_ngat), .B(G2515_553_ngat), .Y(G2524_576_gat) );
AND3XL U_g352 (.A(G1525_540_gat), .B(G1481_543_gat), .C(G1490_542_gat), .Y(G1541_577_gat) );
INVXL U_g353 (.A(G1525_540_gat), .Y(G1528_578_gat) );
INVXL U_g354 (.A(G1521_541_gat), .Y(G1524_579_gat) );
AND3XL U_g355 (.A(G1521_541_gat), .B(G1477_421_gat), .C(G1486_420_gat), .Y(G1538_580_gat) );
AND2XL U_g356 (.A(G553_554_gat), .B(G551_544_gat), .Y(G319_656_gat) );
BUFX20 U_g357 (.A(G1473_545_gat), .Y(G2665_582_gat) );
OR2XL U_g358 (.A(G1473_545_ngat), .B(G2103_247_ngat), .Y(G1218_583_gat) );
INVXL U_g359 (.A(G2730_546_gat), .Y(G2734_584_gat) );
OR2XL U_g360 (.A(G1470_562_ngat), .B(G2099_249_ngat), .Y(G1213_585_gat) );
BUFX20 U_g361 (.A(G1795_547_gat), .Y(G1810_586_gat) );
BUFX20 U_g362 (.A(G1795_547_gat), .Y(G1806_587_gat) );
INVXL U_g363 (.A(G1786_548_gat), .Y(G1790_588_gat) );
INVXL U_g364 (.A(G2525_549_gat), .Y(G2531_589_gat) );
INVXL U_g365 (.A(G2528_550_gat), .Y(G2532_590_gat) );
BUFX20 U_g366 (.A(G1518_551_gat), .Y(G1533_591_gat) );
BUFX20 U_g367 (.A(G1518_551_gat), .Y(G1529_592_gat) );
INVXL U_g368 (.A(G1509_552_gat), .Y(G1513_593_gat) );
AND2XL U_g369 (.A(G1385_283_gat), .B(G1461_559_gat), .Y(G1387_594_gat) );
INVXL U_g370 (.A(G2515_553_gat), .Y(G2521_595_gat) );
AND2XL U_g371 (.A(G875_290_gat), .B(G841_573_gat), .Y(G885_596_gat) );
AND2XL U_g372 (.A(G875_290_gat), .B(G846_565_gat), .Y(G887_597_gat) );
AND2XL U_g373 (.A(G868_198_gat), .B(G1327_568_gat), .Y(G893_598_gat) );
AND2XL U_g374 (.A(G860_197_gat), .B(G841_573_gat), .Y(G152_599_gat) );
AND2XL U_g375 (.A(G860_197_gat), .B(G846_565_gat), .Y(G147_600_gat) );
AND2XL U_g376 (.A(G860_197_gat), .B(G838_564_gat), .Y(G144_601_gat) );
INVXL U_g377 (.A(G2634_555_gat), .Y(G2638_602_gat) );
BUFX20 U_g378 (.A(G1701_556_gat), .Y(G2642_603_gat) );
BUFX20 U_g379 (.A(G1704_557_gat), .Y(G1250_604_gat) );
BUFX20 U_g380 (.A(G1704_557_gat), .Y(G2639_605_gat) );
BUFX20 U_g381 (.A(G1707_558_gat), .Y(G2650_606_gat) );
BUFX20 U_g382 (.A(G1461_559_gat), .Y(G2647_608_gat) );
INVXL U_g383 (.A(G1464_560_gat), .Y(G1389_610_gat) );
BUFX20 U_g384 (.A(G1464_560_gat), .Y(G2658_611_gat) );
BUFX20 U_g385 (.A(G1467_561_gat), .Y(G2655_613_gat) );
BUFX20 U_g386 (.A(G1470_562_gat), .Y(G2668_614_gat) );
BUFX20 U_g387 (.A(G1698_563_gat), .Y(G2631_615_gat) );
BUFX20 U_g388 (.A(G838_564_gat), .Y(G516_616_gat) );
INVXL U_g389 (.A(G838_564_gat), .Y(G1028_617_gat) );
INVXL U_g390 (.A(G846_565_gat), .Y(G1035_618_gat) );
INVXL U_g391 (.A(G846_565_gat), .Y(G852_619_gat) );
BUFX20 U_g392 (.A(G854_566_gat), .Y(G299_692_gat) );
BUFX20 U_g393 (.A(G857_567_gat), .Y(G301_694_gat) );
BUFX20 U_g394 (.A(G1327_568_gat), .Y(G286_696_gat) );
BUFX20 U_g395 (.A(G1329_569_gat), .Y(G303_698_gat) );
BUFX20 U_g396 (.A(G1331_570_gat), .Y(G288_700_gat) );
BUFX20 U_g397 (.A(G1333_571_gat), .Y(G305_702_gat) );
BUFX20 U_g398 (.A(G1335_572_gat), .Y(G290_704_gat) );
INVXL U_g399 (.A(G841_573_gat), .Y(G1031_630_gat) );
BUFX20 U_g400 (.A(G841_573_gat), .Y(G2154_631_gat) );
AND2XL U_g401 (.A(G2012_313_gat), .B(G1467_561_gat), .Y(G2036_632_gat) );
AND2XL U_g402 (.A(G2012_313_gat), .B(G1464_560_gat), .Y(G2034_633_gat) );
AND2XL U_g403 (.A(G2012_313_gat), .B(G1461_559_gat), .Y(G2032_634_gat) );
AND2XL U_g404 (.A(G2012_313_gat), .B(G1470_562_gat), .Y(G2038_635_gat) );
AND2XL U_g405 (.A(G2001_314_gat), .B(G1698_563_gat), .Y(G2024_636_gat) );
AND2XL U_g406 (.A(G2001_314_gat), .B(G1707_558_gat), .Y(G2030_637_gat) );
AND2XL U_g407 (.A(G2001_314_gat), .B(G1704_557_gat), .Y(G2028_638_gat) );
AND2XL U_g408 (.A(G2001_314_gat), .B(G1701_556_gat), .Y(G2026_639_gat) );
AND2XL U_g409 (.A(G1721_315_gat), .B(G1331_570_gat), .Y(G1747_640_gat) );
AND2XL U_g410 (.A(G1721_315_gat), .B(G1329_569_gat), .Y(G1745_641_gat) );
AND2XL U_g411 (.A(G1721_315_gat), .B(G1327_568_gat), .Y(G1743_642_gat) );
AND2XL U_g412 (.A(G1721_315_gat), .B(G1335_572_gat), .Y(G1751_643_gat) );
AND2XL U_g413 (.A(G1721_315_gat), .B(G1333_571_gat), .Y(G1749_644_gat) );
AND2XL U_g414 (.A(G1710_316_gat), .B(G841_573_gat), .Y(G1735_645_gat) );
AND2XL U_g415 (.A(G1710_316_gat), .B(G857_567_gat), .Y(G1741_646_gat) );
AND2XL U_g416 (.A(G1710_316_gat), .B(G854_566_gat), .Y(G1739_647_gat) );
AND2XL U_g417 (.A(G1710_316_gat), .B(G846_565_gat), .Y(G1737_648_gat) );
AND3XL U_g418 (.A(G1806_587_gat), .B(G1777_537_gat), .C(G1786_548_gat), .Y(G1821_649_gat) );
AND3XL U_g419 (.A(G1810_586_gat), .B(G1781_574_gat), .C(G1790_588_gat), .Y(G1824_650_gat) );
AND3XL U_g420 (.A(G1529_592_gat), .B(G1500_538_gat), .C(G1509_552_gat), .Y(G1544_651_gat) );
AND3XL U_g421 (.A(G1533_591_gat), .B(G1504_575_gat), .C(G1513_593_gat), .Y(G1547_652_gat) );
OR2XL U_g422 (.A(G2521_595_ngat), .B(G2518_418_ngat), .Y(G2523_653_gat) );
AND3XL U_g423 (.A(G1524_579_gat), .B(G1486_420_gat), .C(G1481_543_gat), .Y(G1537_654_gat) );
AND3XL U_g424 (.A(G1528_578_gat), .B(G1490_542_gat), .C(G1477_421_gat), .Y(G1540_655_gat) );
AND2XL U_g425 (.A(G1473_545_gat), .B(G1218_583_gat), .Y(G1234_657_gat) );
INVXL U_g426 (.A(G2665_582_gat), .Y(G2671_658_gat) );
AND2XL U_g427 (.A(G1218_583_gat), .B(G2103_247_gat), .Y(G1232_659_gat) );
AND2XL U_g428 (.A(G1213_585_gat), .B(G2099_249_gat), .Y(G1225_660_gat) );
INVXL U_g429 (.A(G1810_586_gat), .Y(G1813_661_gat) );
INVXL U_g430 (.A(G1806_587_gat), .Y(G1809_662_gat) );
OR2XL U_g431 (.A(G2532_590_ngat), .B(G2525_549_ngat), .Y(G2534_663_gat) );
OR2XL U_g432 (.A(G2531_589_ngat), .B(G2528_550_ngat), .Y(G2533_664_gat) );
INVXL U_g433 (.A(G1533_591_gat), .Y(G1536_665_gat) );
INVXL U_g434 (.A(G1529_592_gat), .Y(G1532_666_gat) );
INVXL U_g435 (.A(G1387_594_gat), .Y(G466_667_gat) );
AND2XL U_g436 (.A(G875_290_gat), .B(G516_616_gat), .Y(G883_668_gat) );
AND2XL U_g437 (.A(G875_290_gat), .B(G299_692_gat), .Y(G891_669_gat) );
AND2XL U_g438 (.A(G868_198_gat), .B(G301_694_gat), .Y(G889_670_gat) );
OR2XL U_g439 (.A(G852_619_ngat), .B(G560_295_ngat), .Y(G562_672_gat) );
AND4XL U_g440 (.A(G547_415_gat), .B(G319_656_gat), .C(G483_191_gat), .D(G480_292_gat), .Y(G187_673_gat) );
OR2XL U_g441 (.A(G2638_602_ngat), .B(G2631_615_ngat), .Y(G1753_674_gat) );
INVXL U_g442 (.A(G2642_603_gat), .Y(G2646_675_gat) );
INVXL U_g443 (.A(G2639_605_gat), .Y(G2645_676_gat) );
INVXL U_g444 (.A(G2650_606_gat), .Y(G2654_677_gat) );
INVXL U_g445 (.A(G2647_608_gat), .Y(G2653_678_gat) );
INVXL U_g446 (.A(G2658_611_gat), .Y(G2662_679_gat) );
INVXL U_g447 (.A(G2655_613_gat), .Y(G2661_680_gat) );
AND2XL U_g448 (.A(G1470_562_gat), .B(G1213_585_gat), .Y(G1227_681_gat) );
INVXL U_g449 (.A(G2668_614_gat), .Y(G2672_682_gat) );
INVXL U_g450 (.A(G2631_615_gat), .Y(G2637_683_gat) );
BUFX20 U_g451 (.A(G516_616_gat), .Y(G2235_684_gat) );
BUFX20 U_g452 (.A(G1028_617_gat), .Y(G2110_685_gat) );
BUFX20 U_g453 (.A(G1028_617_gat), .Y(G2164_686_gat) );
BUFX20 U_g454 (.A(G1035_618_gat), .Y(G2350_687_gat) );
BUFX20 U_g455 (.A(G1035_618_gat), .Y(G2118_688_gat) );
BUFX20 U_g456 (.A(G1035_618_gat), .Y(G2262_689_gat) );
BUFX20 U_g457 (.A(G1035_618_gat), .Y(G2172_690_gat) );
INVXL U_g458 (.A(G852_619_gat), .Y(G2151_691_gat) );
INVXL U_g459 (.A(G299_692_gat), .Y(G1043_693_gat) );
INVXL U_g460 (.A(G301_694_gat), .Y(G1051_695_gat) );
INVXL U_g461 (.A(G286_696_gat), .Y(G2123_697_gat) );
INVXL U_g462 (.A(G303_698_gat), .Y(G1062_699_gat) );
INVXL U_g463 (.A(G288_700_gat), .Y(G1068_701_gat) );
INVXL U_g464 (.A(G305_702_gat), .Y(G1074_703_gat) );
INVXL U_g465 (.A(G290_704_gat), .Y(G1080_705_gat) );
BUFX20 U_g466 (.A(G1031_630_gat), .Y(G2107_706_gat) );
BUFX20 U_g467 (.A(G1031_630_gat), .Y(G2161_707_gat) );
INVXL U_g468 (.A(G2154_631_gat), .Y(G2158_708_gat) );
AND3XL U_g469 (.A(G40_29_gat), .B(G1387_594_gat), .C(G1389_610_gat), .Y(G456_709_gat) );
AND4XL U_g470 (.A(G319_656_gat), .B(G36_27_gat), .C(G483_191_gat), .D(G480_292_gat), .Y(G175_710_gat) );
OR2XL U_g471 (.A(G2036_632_gat), .B(G2035_519_gat), .Y(G2778_711_gat) );
OR2XL U_g472 (.A(G2034_633_gat), .B(G2033_520_gat), .Y(G2770_712_gat) );
OR2XL U_g473 (.A(G2030_637_gat), .B(G2029_521_gat), .Y(G2754_713_gat) );
OR2XL U_g474 (.A(G2026_639_gat), .B(G2025_522_gat), .Y(G2738_714_gat) );
OR2XL U_g475 (.A(G2038_635_gat), .B(G2037_523_gat), .Y(G2065_715_gat) );
OR2XL U_g476 (.A(G2032_634_gat), .B(G2031_524_gat), .Y(G2762_716_gat) );
OR2XL U_g477 (.A(G2028_638_gat), .B(G2027_525_gat), .Y(G2746_717_gat) );
OR2XL U_g478 (.A(G2024_636_gat), .B(G2023_526_gat), .Y(G2626_718_gat) );
OR2XL U_g479 (.A(G1751_643_gat), .B(G1750_527_gat), .Y(G2618_719_gat) );
OR2XL U_g480 (.A(G1747_640_gat), .B(G1746_528_gat), .Y(G2602_720_gat) );
OR2XL U_g481 (.A(G1745_641_gat), .B(G1744_529_gat), .Y(G2594_721_gat) );
OR2XL U_g482 (.A(G1743_642_gat), .B(G1742_530_gat), .Y(G2586_722_gat) );
OR2XL U_g483 (.A(G1739_647_gat), .B(G1738_531_gat), .Y(G2570_723_gat) );
OR2XL U_g484 (.A(G1735_645_gat), .B(G1734_532_gat), .Y(G2554_724_gat) );
OR2XL U_g485 (.A(G1749_644_gat), .B(G1748_534_gat), .Y(G2610_725_gat) );
OR2XL U_g486 (.A(G1741_646_gat), .B(G1740_535_gat), .Y(G2578_726_gat) );
OR2XL U_g487 (.A(G1737_648_gat), .B(G1736_536_gat), .Y(G2562_727_gat) );
AND3XL U_g488 (.A(G1813_661_gat), .B(G1790_588_gat), .C(G1777_537_gat), .Y(G1823_728_gat) );
AND3XL U_g489 (.A(G1536_665_gat), .B(G1513_593_gat), .C(G1500_538_gat), .Y(G1546_729_gat) );
OR2XL U_g490 (.A(G2524_576_ngat), .B(G2523_653_ngat), .Y(G2538_730_gat) );
AND2XL U_g491 (.A(G1541_577_ngat), .B(G1540_655_ngat), .Y(G1542_731_gat) );
AND2XL U_g492 (.A(G1538_580_ngat), .B(G1537_654_ngat), .Y(G1539_732_gat) );
OR2XL U_g493 (.A(G1234_657_gat), .B(G1232_659_gat), .Y(G1235_733_gat) );
OR2XL U_g494 (.A(G2672_682_ngat), .B(G2665_582_ngat), .Y(G2674_734_gat) );
OR2XL U_g495 (.A(G1227_681_gat), .B(G1225_660_gat), .Y(G1228_735_gat) );
OR2XL U_g496 (.A(G2781_429_ngat), .B(G2778_711_ngat), .Y(G2059_736_gat) );
OR2XL U_g497 (.A(G2773_431_ngat), .B(G2770_712_ngat), .Y(G2055_737_gat) );
OR2XL U_g498 (.A(G2765_433_ngat), .B(G2762_716_ngat), .Y(G2051_738_gat) );
AND3XL U_g499 (.A(G1809_662_gat), .B(G1786_548_gat), .C(G1781_574_gat), .Y(G1820_739_gat) );
OR2XL U_g500 (.A(G2757_435_ngat), .B(G2754_713_ngat), .Y(G2047_740_gat) );
OR2XL U_g501 (.A(G2749_437_ngat), .B(G2746_717_ngat), .Y(G2043_741_gat) );
OR2XL U_g502 (.A(G2741_438_ngat), .B(G2738_714_ngat), .Y(G2039_742_gat) );
OR2XL U_g503 (.A(G2534_663_ngat), .B(G2533_664_ngat), .Y(G2546_743_gat) );
OR2XL U_g504 (.A(G2629_440_ngat), .B(G2626_718_ngat), .Y(G1597_744_gat) );
OR2XL U_g505 (.A(G2621_442_ngat), .B(G2618_719_ngat), .Y(G1593_745_gat) );
OR2XL U_g506 (.A(G2613_444_ngat), .B(G2610_725_ngat), .Y(G1589_746_gat) );
OR2XL U_g507 (.A(G2605_446_ngat), .B(G2602_720_ngat), .Y(G1585_747_gat) );
OR2XL U_g508 (.A(G2597_448_ngat), .B(G2594_721_ngat), .Y(G1581_748_gat) );
OR2XL U_g509 (.A(G2589_450_ngat), .B(G2586_722_ngat), .Y(G1577_749_gat) );
AND3XL U_g510 (.A(G1532_666_gat), .B(G1509_552_gat), .C(G1504_575_gat), .Y(G1543_750_gat) );
OR2XL U_g511 (.A(G2581_452_ngat), .B(G2578_726_ngat), .Y(G1573_751_gat) );
OR2XL U_g512 (.A(G2573_454_ngat), .B(G2570_723_ngat), .Y(G1569_752_gat) );
OR2XL U_g513 (.A(G2565_455_ngat), .B(G2562_727_ngat), .Y(G1565_753_gat) );
OR2XL U_g514 (.A(G2557_457_ngat), .B(G2554_724_ngat), .Y(G1561_754_gat) );
OR2XL U_g515 (.A(G889_670_gat), .B(G887_597_gat), .Y(G897_755_gat) );
OR2XL U_g516 (.A(G893_598_gat), .B(G891_669_gat), .Y(G898_756_gat) );
AND2XL U_g517 (.A(G868_198_gat), .B(G562_672_gat), .Y(G886_757_gat) );
AND2XL U_g518 (.A(G865_291_gat), .B(G562_672_gat), .Y(G146_758_gat) );
INVXL U_g519 (.A(G562_672_gat), .Y(G2207_759_gat) );
BUFX20 U_g520 (.A(G562_672_gat), .Y(G592_760_gat) );
OR2XL U_g521 (.A(G2637_683_ngat), .B(G2634_555_ngat), .Y(G1752_762_gat) );
OR2XL U_g522 (.A(G2645_676_ngat), .B(G2642_603_ngat), .Y(G1761_763_gat) );
OR2XL U_g523 (.A(G2646_675_ngat), .B(G2639_605_ngat), .Y(G1762_764_gat) );
OR2XL U_g524 (.A(G2653_678_ngat), .B(G2650_606_ngat), .Y(G1770_765_gat) );
OR2XL U_g525 (.A(G2654_677_ngat), .B(G2647_608_ngat), .Y(G1771_766_gat) );
OR2XL U_g526 (.A(G2661_680_ngat), .B(G2658_611_ngat), .Y(G2663_767_gat) );
OR2XL U_g527 (.A(G2662_679_ngat), .B(G2655_613_ngat), .Y(G2664_768_gat) );
OR2XL U_g528 (.A(G2671_658_ngat), .B(G2668_614_ngat), .Y(G2673_769_gat) );
INVXL U_g529 (.A(G2235_684_gat), .Y(G2241_770_gat) );
INVXL U_g530 (.A(G2110_685_gat), .Y(G2114_771_gat) );
INVXL U_g531 (.A(G2164_686_gat), .Y(G2168_772_gat) );
INVXL U_g532 (.A(G2350_687_gat), .Y(G2354_773_gat) );
INVXL U_g533 (.A(G2118_688_gat), .Y(G2122_774_gat) );
INVXL U_g534 (.A(G2262_689_gat), .Y(G2266_775_gat) );
INVXL U_g535 (.A(G2172_690_gat), .Y(G2176_776_gat) );
INVXL U_g536 (.A(G2151_691_gat), .Y(G2157_777_gat) );
OR2XL U_g537 (.A(G2158_708_ngat), .B(G2151_691_ngat), .Y(G2160_778_gat) );
BUFX20 U_g538 (.A(G1043_693_gat), .Y(G2342_779_gat) );
BUFX20 U_g539 (.A(G1043_693_gat), .Y(G2115_780_gat) );
BUFX20 U_g540 (.A(G1043_693_gat), .Y(G2254_781_gat) );
BUFX20 U_g541 (.A(G1043_693_gat), .Y(G2169_782_gat) );
BUFX20 U_g542 (.A(G1051_695_gat), .Y(G2422_783_gat) );
BUFX20 U_g543 (.A(G1051_695_gat), .Y(G2334_784_gat) );
BUFX20 U_g544 (.A(G1051_695_gat), .Y(G2126_785_gat) );
INVXL U_g545 (.A(G2123_697_gat), .Y(G2129_786_gat) );
BUFX20 U_g546 (.A(G1062_699_gat), .Y(G2134_787_gat) );
BUFX20 U_g547 (.A(G1062_699_gat), .Y(G2180_788_gat) );
BUFX20 U_g548 (.A(G1068_701_gat), .Y(G2131_789_gat) );
BUFX20 U_g549 (.A(G1068_701_gat), .Y(G2177_790_gat) );
BUFX20 U_g550 (.A(G1074_703_gat), .Y(G2144_791_gat) );
BUFX20 U_g551 (.A(G1074_703_gat), .Y(G2190_792_gat) );
BUFX20 U_g552 (.A(G1080_705_gat), .Y(G2141_793_gat) );
BUFX20 U_g553 (.A(G1080_705_gat), .Y(G2187_794_gat) );
INVXL U_g554 (.A(G2107_706_gat), .Y(G2113_795_gat) );
INVXL U_g555 (.A(G2161_707_gat), .Y(G2167_796_gat) );
AND3XL U_g556 (.A(G466_667_gat), .B(G1389_610_gat), .C(G40_29_gat), .Y(G468_797_gat) );
BUFX20 U_g557 (.A(G456_709_gat), .Y(G995_798_gat) );
INVXL U_g558 (.A(G456_709_gat), .Y(G1006_799_gat) );
INVXL U_g559 (.A(G456_709_gat), .Y(G743_800_gat) );
BUFX20 U_g560 (.A(G456_709_gat), .Y(G749_801_gat) );
INVXL U_g561 (.A(G456_709_gat), .Y(G462_802_gat) );
INVXL U_g562 (.A(G2778_711_gat), .Y(G2782_804_gat) );
INVXL U_g563 (.A(G2770_712_gat), .Y(G2774_805_gat) );
INVXL U_g564 (.A(G2754_713_gat), .Y(G2758_806_gat) );
INVXL U_g565 (.A(G2738_714_gat), .Y(G2742_807_gat) );
INVXL U_g566 (.A(G2762_716_gat), .Y(G2766_808_gat) );
INVXL U_g567 (.A(G2746_717_gat), .Y(G2750_809_gat) );
INVXL U_g568 (.A(G2626_718_gat), .Y(G2630_810_gat) );
INVXL U_g569 (.A(G2618_719_gat), .Y(G2622_811_gat) );
INVXL U_g570 (.A(G2602_720_gat), .Y(G2606_812_gat) );
INVXL U_g571 (.A(G2594_721_gat), .Y(G2598_813_gat) );
INVXL U_g572 (.A(G2586_722_gat), .Y(G2590_814_gat) );
INVXL U_g573 (.A(G2570_723_gat), .Y(G2574_815_gat) );
INVXL U_g574 (.A(G2554_724_gat), .Y(G2558_816_gat) );
INVXL U_g575 (.A(G2610_725_gat), .Y(G2614_817_gat) );
INVXL U_g576 (.A(G2578_726_gat), .Y(G2582_818_gat) );
INVXL U_g577 (.A(G2562_727_gat), .Y(G2566_819_gat) );
AND2XL U_g578 (.A(G1821_649_ngat), .B(G1820_739_ngat), .Y(G1822_820_gat) );
AND2XL U_g579 (.A(G1824_650_ngat), .B(G1823_728_ngat), .Y(G1825_821_gat) );
AND2XL U_g580 (.A(G1544_651_ngat), .B(G1543_750_ngat), .Y(G1545_822_gat) );
AND2XL U_g581 (.A(G1547_652_ngat), .B(G1546_729_ngat), .Y(G1548_823_gat) );
INVXL U_g582 (.A(G2538_730_gat), .Y(G2542_824_gat) );
OR2XL U_g583 (.A(G1539_732_ngat), .B(G1542_731_ngat), .Y(G2535_825_gat) );
INVXL U_g584 (.A(G1235_733_gat), .Y(G1245_826_gat) );
OR2XL U_g585 (.A(G2674_734_ngat), .B(G2673_769_ngat), .Y(G2709_827_gat) );
INVXL U_g586 (.A(G1228_735_gat), .Y(G1243_828_gat) );
OR2XL U_g587 (.A(G2782_804_ngat), .B(G2775_341_ngat), .Y(G2060_829_gat) );
OR2XL U_g588 (.A(G2774_805_ngat), .B(G2767_343_ngat), .Y(G2056_830_gat) );
OR2XL U_g589 (.A(G2766_808_ngat), .B(G2759_345_ngat), .Y(G2052_831_gat) );
OR2XL U_g590 (.A(G2758_806_ngat), .B(G2751_347_ngat), .Y(G2048_832_gat) );
OR2XL U_g591 (.A(G2750_809_ngat), .B(G2743_350_ngat), .Y(G2044_833_gat) );
OR2XL U_g592 (.A(G2742_807_ngat), .B(G2735_352_ngat), .Y(G2040_834_gat) );
INVXL U_g593 (.A(G2546_743_gat), .Y(G2550_835_gat) );
OR2XL U_g594 (.A(G2630_810_ngat), .B(G2623_354_ngat), .Y(G1598_836_gat) );
OR2XL U_g595 (.A(G2622_811_ngat), .B(G2615_356_ngat), .Y(G1594_837_gat) );
OR2XL U_g596 (.A(G2614_817_ngat), .B(G2607_358_ngat), .Y(G1590_838_gat) );
OR2XL U_g597 (.A(G2606_812_ngat), .B(G2599_360_ngat), .Y(G1586_839_gat) );
OR2XL U_g598 (.A(G2598_813_ngat), .B(G2591_362_ngat), .Y(G1582_840_gat) );
OR2XL U_g599 (.A(G2590_814_ngat), .B(G2583_364_ngat), .Y(G1578_841_gat) );
OR2XL U_g600 (.A(G2582_818_ngat), .B(G2575_366_ngat), .Y(G1574_842_gat) );
OR2XL U_g601 (.A(G2574_815_ngat), .B(G2567_368_ngat), .Y(G1570_843_gat) );
OR2XL U_g602 (.A(G2566_819_ngat), .B(G2559_370_ngat), .Y(G1566_844_gat) );
OR2XL U_g603 (.A(G2558_816_ngat), .B(G2551_372_ngat), .Y(G1562_845_gat) );
OR2XL U_g604 (.A(G886_757_gat), .B(G885_596_gat), .Y(G896_846_gat) );
INVXL U_g605 (.A(G2207_759_gat), .Y(G2213_852_gat) );
INVXL U_g606 (.A(G592_760_gat), .Y(G596_853_gat) );
OR2XL U_g607 (.A(G1753_674_ngat), .B(G1752_762_ngat), .Y(G1754_854_gat) );
AND2XL U_g608 (.A(G743_800_gat), .B(G1701_556_gat), .Y(G502_855_gat) );
AND2XL U_g609 (.A(G1006_799_gat), .B(G1701_556_gat), .Y(G729_856_gat) );
OR2XL U_g610 (.A(G1762_764_ngat), .B(G1761_763_ngat), .Y(G1763_857_gat) );
AND2XL U_g611 (.A(G743_800_gat), .B(G1250_604_gat), .Y(G508_858_gat) );
AND2XL U_g612 (.A(G1006_799_gat), .B(G1250_604_gat), .Y(G735_859_gat) );
OR2XL U_g613 (.A(G1771_766_ngat), .B(G1770_765_ngat), .Y(G1772_860_gat) );
OR2XL U_g614 (.A(G2664_768_ngat), .B(G2663_767_ngat), .Y(G2712_861_gat) );
AND2XL U_g615 (.A(G743_800_gat), .B(G1698_563_gat), .Y(G496_862_gat) );
AND2XL U_g616 (.A(G1006_799_gat), .B(G1698_563_gat), .Y(G723_863_gat) );
OR2XL U_g617 (.A(G2113_795_ngat), .B(G2110_685_ngat), .Y(G569_864_gat) );
OR2XL U_g618 (.A(G2167_796_ngat), .B(G2164_686_ngat), .Y(G599_865_gat) );
OR2XL U_g619 (.A(G2122_774_ngat), .B(G2115_780_ngat), .Y(G579_866_gat) );
OR2XL U_g620 (.A(G2176_776_ngat), .B(G2169_782_ngat), .Y(G609_867_gat) );
INVXL U_g621 (.A(G2342_779_gat), .Y(G2346_868_gat) );
INVXL U_g622 (.A(G2115_780_gat), .Y(G2121_869_gat) );
INVXL U_g623 (.A(G2254_781_gat), .Y(G2258_870_gat) );
INVXL U_g624 (.A(G2169_782_gat), .Y(G2175_871_gat) );
INVXL U_g625 (.A(G2422_783_gat), .Y(G2426_872_gat) );
INVXL U_g626 (.A(G2334_784_gat), .Y(G2338_873_gat) );
OR2XL U_g627 (.A(G2129_786_ngat), .B(G2126_785_ngat), .Y(G587_874_gat) );
INVXL U_g628 (.A(G2126_785_gat), .Y(G2130_875_gat) );
AND2XL U_g629 (.A(G749_801_gat), .B(G286_696_gat), .Y(G765_876_gat) );
AND2XL U_g630 (.A(G995_798_gat), .B(G286_696_gat), .Y(G1014_877_gat) );
AND2XL U_g631 (.A(G749_801_gat), .B(G303_698_gat), .Y(G769_878_gat) );
AND2XL U_g632 (.A(G995_798_gat), .B(G303_698_gat), .Y(G1018_879_gat) );
INVXL U_g633 (.A(G2134_787_gat), .Y(G2138_880_gat) );
INVXL U_g634 (.A(G2180_788_gat), .Y(G2184_881_gat) );
INVXL U_g635 (.A(G2131_789_gat), .Y(G2137_882_gat) );
INVXL U_g636 (.A(G2177_790_gat), .Y(G2183_883_gat) );
INVXL U_g637 (.A(G2144_791_gat), .Y(G2148_884_gat) );
INVXL U_g638 (.A(G2190_792_gat), .Y(G2194_885_gat) );
AND2XL U_g639 (.A(G743_800_gat), .B(G290_704_gat), .Y(G490_886_gat) );
AND2XL U_g640 (.A(G1006_799_gat), .B(G290_704_gat), .Y(G717_887_gat) );
INVXL U_g641 (.A(G2141_793_gat), .Y(G2147_888_gat) );
INVXL U_g642 (.A(G2187_794_gat), .Y(G2193_889_gat) );
OR2XL U_g643 (.A(G2114_771_ngat), .B(G2107_706_ngat), .Y(G570_890_gat) );
OR2XL U_g644 (.A(G2168_772_ngat), .B(G2161_707_ngat), .Y(G600_891_gat) );
OR2XL U_g645 (.A(G2157_777_ngat), .B(G2154_631_ngat), .Y(G2159_892_gat) );
BUFX20 U_g646 (.A(G468_797_gat), .Y(G1257_893_gat) );
BUFX20 U_g647 (.A(G468_797_gat), .Y(G1258_894_gat) );
INVXL U_g648 (.A(G995_798_gat), .Y(G999_895_gat) );
INVXL U_g649 (.A(G749_801_gat), .Y(G753_896_gat) );
BUFX20 U_g650 (.A(G462_802_gat), .Y(G475_897_gat) );
BUFX20 U_g651 (.A(G462_802_gat), .Y(G1337_898_gat) );
OR2XL U_g652 (.A(G1822_820_ngat), .B(G1825_821_ngat), .Y(G2727_899_gat) );
OR2XL U_g653 (.A(G1545_822_ngat), .B(G1548_823_ngat), .Y(G2543_900_gat) );
OR2XL U_g654 (.A(G2542_824_ngat), .B(G2535_825_ngat), .Y(G1550_901_gat) );
INVXL U_g655 (.A(G2535_825_gat), .Y(G2541_902_gat) );
AND2XL U_g656 (.A(G1245_826_gat), .B(G1235_733_gat), .Y(G1094_903_gat) );
INVXL U_g657 (.A(G2709_827_gat), .Y(G2715_904_gat) );
AND2XL U_g658 (.A(G1243_828_gat), .B(G1228_735_gat), .Y(G1096_905_gat) );
OR2XL U_g659 (.A(G2060_829_ngat), .B(G2059_736_ngat), .Y(G2061_906_gat) );
OR2XL U_g660 (.A(G2056_830_ngat), .B(G2055_737_ngat), .Y(G2057_907_gat) );
OR2XL U_g661 (.A(G2052_831_ngat), .B(G2051_738_ngat), .Y(G2053_908_gat) );
OR2XL U_g662 (.A(G2048_832_ngat), .B(G2047_740_ngat), .Y(G2049_909_gat) );
OR2XL U_g663 (.A(G2044_833_ngat), .B(G2043_741_ngat), .Y(G2045_910_gat) );
OR2XL U_g664 (.A(G2040_834_ngat), .B(G2039_742_ngat), .Y(G2041_911_gat) );
OR2XL U_g665 (.A(G1598_836_ngat), .B(G1597_744_ngat), .Y(G1599_912_gat) );
OR2XL U_g666 (.A(G1594_837_ngat), .B(G1593_745_ngat), .Y(G1595_913_gat) );
OR2XL U_g667 (.A(G1590_838_ngat), .B(G1589_746_ngat), .Y(G1591_914_gat) );
OR2XL U_g668 (.A(G1586_839_ngat), .B(G1585_747_ngat), .Y(G1587_915_gat) );
OR2XL U_g669 (.A(G1582_840_ngat), .B(G1581_748_ngat), .Y(G1583_916_gat) );
OR2XL U_g670 (.A(G1578_841_ngat), .B(G1577_749_ngat), .Y(G1579_917_gat) );
OR2XL U_g671 (.A(G1574_842_ngat), .B(G1573_751_ngat), .Y(G1575_918_gat) );
OR2XL U_g672 (.A(G1570_843_ngat), .B(G1569_752_ngat), .Y(G1571_919_gat) );
OR2XL U_g673 (.A(G1566_844_ngat), .B(G1565_753_ngat), .Y(G1567_920_gat) );
OR2XL U_g674 (.A(G1562_845_ngat), .B(G1561_754_ngat), .Y(G1563_921_gat) );
INVXL U_g675 (.A(G1754_854_gat), .Y(G1758_924_gat) );
INVXL U_g676 (.A(G1763_857_gat), .Y(G1767_925_gat) );
BUFX20 U_g677 (.A(G1772_860_gat), .Y(G1802_926_gat) );
BUFX20 U_g678 (.A(G1772_860_gat), .Y(G1798_927_gat) );
INVXL U_g679 (.A(G2712_861_gat), .Y(G2716_928_gat) );
OR2XL U_g680 (.A(G570_890_ngat), .B(G569_864_ngat), .Y(G571_929_gat) );
OR2XL U_g681 (.A(G600_891_ngat), .B(G599_865_ngat), .Y(G601_930_gat) );
OR2XL U_g682 (.A(G2121_869_ngat), .B(G2118_688_ngat), .Y(G578_931_gat) );
OR2XL U_g683 (.A(G2175_871_ngat), .B(G2172_690_ngat), .Y(G608_932_gat) );
OR2XL U_g684 (.A(G2160_778_ngat), .B(G2159_892_ngat), .Y(G2210_933_gat) );
AND2XL U_g685 (.A(G753_896_gat), .B(G286_696_gat), .Y(G763_934_gat) );
AND2XL U_g686 (.A(G999_895_gat), .B(G286_696_gat), .Y(G1012_935_gat) );
OR2XL U_g687 (.A(G2130_875_ngat), .B(G2123_697_ngat), .Y(G588_936_gat) );
AND2XL U_g688 (.A(G753_896_gat), .B(G303_698_gat), .Y(G767_937_gat) );
AND2XL U_g689 (.A(G999_895_gat), .B(G303_698_gat), .Y(G1016_938_gat) );
OR2XL U_g690 (.A(G2137_882_ngat), .B(G2134_787_ngat), .Y(G2139_939_gat) );
OR2XL U_g691 (.A(G2183_883_ngat), .B(G2180_788_ngat), .Y(G2185_940_gat) );
AND2XL U_g692 (.A(G753_896_gat), .B(G288_700_gat), .Y(G531_941_gat) );
AND2XL U_g693 (.A(G999_895_gat), .B(G288_700_gat), .Y(G705_942_gat) );
OR2XL U_g694 (.A(G2138_880_ngat), .B(G2131_789_ngat), .Y(G2140_943_gat) );
OR2XL U_g695 (.A(G2184_881_ngat), .B(G2177_790_ngat), .Y(G2186_944_gat) );
AND2XL U_g696 (.A(G753_896_gat), .B(G305_702_gat), .Y(G537_945_gat) );
AND2XL U_g697 (.A(G999_895_gat), .B(G305_702_gat), .Y(G711_946_gat) );
OR2XL U_g698 (.A(G2147_888_ngat), .B(G2144_791_ngat), .Y(G2149_947_gat) );
OR2XL U_g699 (.A(G2193_889_ngat), .B(G2190_792_ngat), .Y(G2195_948_gat) );
OR2XL U_g700 (.A(G2148_884_ngat), .B(G2141_793_ngat), .Y(G2150_949_gat) );
OR2XL U_g701 (.A(G2194_885_ngat), .B(G2187_794_ngat), .Y(G2196_950_gat) );
BUFX20 U_g702 (.A(G1257_893_gat), .Y(G742_951_gat) );
BUFX20 U_g703 (.A(G1257_893_gat), .Y(G1005_952_gat) );
BUFX20 U_g704 (.A(G1258_894_gat), .Y(G1845_953_gat) );
BUFX20 U_g705 (.A(G1258_894_gat), .Y(G1907_954_gat) );
BUFX20 U_g706 (.A(G475_897_gat), .Y(G1836_955_gat) );
BUFX20 U_g707 (.A(G475_897_gat), .Y(G1850_956_gat) );
BUFX20 U_g708 (.A(G475_897_gat), .Y(G1355_957_gat) );
BUFX20 U_g709 (.A(G1337_898_gat), .Y(G1898_958_gat) );
BUFX20 U_g710 (.A(G1337_898_gat), .Y(G1912_959_gat) );
BUFX20 U_g711 (.A(G1337_898_gat), .Y(G1601_960_gat) );
INVXL U_g712 (.A(G2727_899_gat), .Y(G2733_961_gat) );
INVXL U_g713 (.A(G2543_900_gat), .Y(G2549_962_gat) );
OR2XL U_g714 (.A(G2541_902_ngat), .B(G2538_730_ngat), .Y(G1549_963_gat) );
OR2XL U_g715 (.A(G1245_826_gat), .B(G1094_903_gat), .Y(G154_964_gat) );
OR2XL U_g716 (.A(G2716_928_ngat), .B(G2709_827_ngat), .Y(G2718_965_gat) );
OR2XL U_g717 (.A(G2734_584_ngat), .B(G2727_899_ngat), .Y(G1829_966_gat) );
OR2XL U_g718 (.A(G1243_828_gat), .B(G1096_905_gat), .Y(G155_967_gat) );
INVXL U_g719 (.A(G2061_906_gat), .Y(G2062_968_gat) );
INVXL U_g720 (.A(G2057_907_gat), .Y(G2058_969_gat) );
INVXL U_g721 (.A(G2053_908_gat), .Y(G2054_970_gat) );
INVXL U_g722 (.A(G2049_909_gat), .Y(G2050_971_gat) );
AND2XL U_g723 (.A(G1850_956_gat), .B(G2070_260_gat), .Y(G1876_972_gat) );
AND2XL U_g724 (.A(G1912_959_gat), .B(G2070_260_gat), .Y(G1938_973_gat) );
INVXL U_g725 (.A(G2045_910_gat), .Y(G2046_974_gat) );
AND2XL U_g726 (.A(G1850_956_gat), .B(G1999_265_gat), .Y(G1874_975_gat) );
AND2XL U_g727 (.A(G1912_959_gat), .B(G1999_265_gat), .Y(G1936_976_gat) );
INVXL U_g728 (.A(G2041_911_gat), .Y(G2042_977_gat) );
OR2XL U_g729 (.A(G2550_835_ngat), .B(G2543_900_ngat), .Y(G1552_978_gat) );
AND2XL U_g730 (.A(G1850_956_gat), .B(G1994_267_gat), .Y(G1872_979_gat) );
AND2XL U_g731 (.A(G1912_959_gat), .B(G1994_267_gat), .Y(G1934_980_gat) );
INVXL U_g732 (.A(G1599_912_gat), .Y(G1600_981_gat) );
AND2XL U_g733 (.A(G1850_956_gat), .B(G1989_269_gat), .Y(G1870_982_gat) );
AND2XL U_g734 (.A(G1912_959_gat), .B(G1989_269_gat), .Y(G1932_983_gat) );
INVXL U_g735 (.A(G1595_913_gat), .Y(G1596_984_gat) );
AND2XL U_g736 (.A(G1836_955_gat), .B(G1984_271_gat), .Y(G1868_985_gat) );
AND2XL U_g737 (.A(G1898_958_gat), .B(G1984_271_gat), .Y(G1930_986_gat) );
INVXL U_g738 (.A(G1591_914_gat), .Y(G1592_987_gat) );
AND2XL U_g739 (.A(G1836_955_gat), .B(G1979_273_gat), .Y(G1866_988_gat) );
AND2XL U_g740 (.A(G1898_958_gat), .B(G1979_273_gat), .Y(G1928_989_gat) );
INVXL U_g741 (.A(G1587_915_gat), .Y(G1588_990_gat) );
AND2XL U_g742 (.A(G1836_955_gat), .B(G1974_275_gat), .Y(G1863_991_gat) );
AND2XL U_g743 (.A(G1898_958_gat), .B(G1974_275_gat), .Y(G1925_992_gat) );
INVXL U_g744 (.A(G1583_916_gat), .Y(G1584_993_gat) );
AND2XL U_g745 (.A(G1836_955_gat), .B(G1969_277_gat), .Y(G1858_994_gat) );
AND2XL U_g746 (.A(G1898_958_gat), .B(G1969_277_gat), .Y(G1920_995_gat) );
INVXL U_g747 (.A(G1579_917_gat), .Y(G1580_996_gat) );
AND2XL U_g748 (.A(G1355_957_gat), .B(G1964_279_gat), .Y(G1377_997_gat) );
AND2XL U_g749 (.A(G1601_960_gat), .B(G1964_279_gat), .Y(G1623_998_gat) );
INVXL U_g750 (.A(G1575_918_gat), .Y(G1576_999_gat) );
AND2XL U_g751 (.A(G1355_957_gat), .B(G1959_281_gat), .Y(G1373_1000_gat) );
AND2XL U_g752 (.A(G1601_960_gat), .B(G1959_281_gat), .Y(G1619_1001_gat) );
INVXL U_g753 (.A(G1571_919_gat), .Y(G1572_1002_gat) );
AND2XL U_g754 (.A(G1601_960_gat), .B(G1351_284_gat), .Y(G1615_1003_gat) );
AND2XL U_g755 (.A(G1355_957_gat), .B(G1351_284_gat), .Y(G1369_1004_gat) );
INVXL U_g756 (.A(G1567_920_gat), .Y(G1568_1005_gat) );
AND2XL U_g757 (.A(G1355_957_gat), .B(G1344_286_gat), .Y(G676_1006_gat) );
AND2XL U_g758 (.A(G1601_960_gat), .B(G1344_286_gat), .Y(G1108_1007_gat) );
INVXL U_g759 (.A(G1563_921_gat), .Y(G1564_1008_gat) );
OR2XL U_g760 (.A(G2213_852_ngat), .B(G2210_933_ngat), .Y(G2215_1009_gat) );
AND3XL U_g761 (.A(G1798_927_gat), .B(G1754_854_gat), .C(G1763_857_gat), .Y(G1815_1010_gat) );
AND3XL U_g762 (.A(G1802_926_gat), .B(G1758_924_gat), .C(G1767_925_gat), .Y(G1818_1011_gat) );
AND2XL U_g763 (.A(G742_951_gat), .B(G502_855_gat), .Y(G504_1012_gat) );
AND2XL U_g764 (.A(G1005_952_gat), .B(G729_856_gat), .Y(G731_1013_gat) );
AND2XL U_g765 (.A(G742_951_gat), .B(G508_858_gat), .Y(G510_1014_gat) );
AND2XL U_g766 (.A(G1005_952_gat), .B(G735_859_gat), .Y(G737_1015_gat) );
INVXL U_g767 (.A(G1802_926_gat), .Y(G1805_1016_gat) );
INVXL U_g768 (.A(G1798_927_gat), .Y(G1801_1017_gat) );
OR2XL U_g769 (.A(G2715_904_ngat), .B(G2712_861_ngat), .Y(G2717_1018_gat) );
AND2XL U_g770 (.A(G742_951_gat), .B(G496_862_gat), .Y(G498_1019_gat) );
AND2XL U_g771 (.A(G1005_952_gat), .B(G723_863_gat), .Y(G725_1020_gat) );
INVXL U_g772 (.A(G571_929_gat), .Y(G575_1021_gat) );
INVXL U_g773 (.A(G601_930_gat), .Y(G605_1022_gat) );
OR2XL U_g774 (.A(G579_866_ngat), .B(G578_931_ngat), .Y(G580_1023_gat) );
OR2XL U_g775 (.A(G609_867_ngat), .B(G608_932_ngat), .Y(G610_1024_gat) );
INVXL U_g776 (.A(G2210_933_gat), .Y(G2214_1025_gat) );
OR2XL U_g777 (.A(G588_936_ngat), .B(G587_874_ngat), .Y(G589_1026_gat) );
OR2XL U_g778 (.A(G765_876_gat), .B(G763_934_gat), .Y(G519_1027_gat) );
OR2XL U_g779 (.A(G1014_877_gat), .B(G1012_935_gat), .Y(G693_1028_gat) );
OR2XL U_g780 (.A(G769_878_gat), .B(G767_937_gat), .Y(G525_1029_gat) );
OR2XL U_g781 (.A(G1018_879_gat), .B(G1016_938_gat), .Y(G699_1030_gat) );
OR2XL U_g782 (.A(G2140_943_ngat), .B(G2139_939_ngat), .Y(G2200_1031_gat) );
OR2XL U_g783 (.A(G2186_944_ngat), .B(G2185_940_ngat), .Y(G2220_1032_gat) );
OR2XL U_g784 (.A(G2150_949_ngat), .B(G2149_947_ngat), .Y(G2197_1033_gat) );
OR2XL U_g785 (.A(G2196_950_ngat), .B(G2195_948_ngat), .Y(G2217_1034_gat) );
AND2XL U_g786 (.A(G742_951_gat), .B(G490_886_gat), .Y(G492_1035_gat) );
AND2XL U_g787 (.A(G1005_952_gat), .B(G717_887_gat), .Y(G719_1036_gat) );
INVXL U_g788 (.A(G1836_955_gat), .Y(G1842_1037_gat) );
INVXL U_g789 (.A(G1355_957_gat), .Y(G1361_1038_gat) );
INVXL U_g790 (.A(G1898_958_gat), .Y(G1904_1039_gat) );
INVXL U_g791 (.A(G1601_960_gat), .Y(G1607_1040_gat) );
AND2XL U_g792 (.A(G748_411_gat), .B(G531_941_gat), .Y(G533_1041_gat) );
AND2XL U_g793 (.A(G748_411_gat), .B(G537_945_gat), .Y(G539_1042_gat) );
AND2XL U_g794 (.A(G994_412_gat), .B(G705_942_gat), .Y(G707_1043_gat) );
AND2XL U_g795 (.A(G994_412_gat), .B(G711_946_gat), .Y(G713_1044_gat) );
OR2XL U_g796 (.A(G1550_901_ngat), .B(G1549_963_ngat), .Y(G1091_1045_gat) );
OR2XL U_g797 (.A(G2718_965_ngat), .B(G2717_1018_ngat), .Y(G2722_1047_gat) );
OR2XL U_g798 (.A(G2733_961_ngat), .B(G2730_546_ngat), .Y(G1828_1048_gat) );
AND2XL U_g799 (.A(G1842_1037_gat), .B(G2094_251_gat), .Y(G1861_1049_gat) );
AND2XL U_g800 (.A(G1904_1039_gat), .B(G2094_251_gat), .Y(G1923_1050_gat) );
AND2XL U_g801 (.A(G1842_1037_gat), .B(G2088_253_gat), .Y(G1856_1051_gat) );
AND2XL U_g802 (.A(G1904_1039_gat), .B(G2088_253_gat), .Y(G1918_1052_gat) );
AND5XL U_g803 (.A(G2042_977_gat), .B(G2046_974_gat), .C(G2050_971_gat), .D(G2054_970_gat), .E(G2058_969_gat), .Y(G1558_1053_gat) );
AND2XL U_g804 (.A(G1361_1038_gat), .B(G2082_255_gat), .Y(G1375_1054_gat) );
AND2XL U_g805 (.A(G1607_1040_gat), .B(G2082_255_gat), .Y(G1621_1055_gat) );
AND2XL U_g806 (.A(G1361_1038_gat), .B(G2076_257_gat), .Y(G1371_1056_gat) );
AND2XL U_g807 (.A(G1607_1040_gat), .B(G2076_257_gat), .Y(G1617_1057_gat) );
AND2XL U_g808 (.A(G1361_1038_gat), .B(G2070_260_gat), .Y(G1368_1058_gat) );
AND2XL U_g809 (.A(G1607_1040_gat), .B(G2070_260_gat), .Y(G1614_1059_gat) );
AND2XL U_g810 (.A(G1361_1038_gat), .B(G1999_265_gat), .Y(G675_1060_gat) );
AND2XL U_g811 (.A(G1607_1040_gat), .B(G1999_265_gat), .Y(G1107_1061_gat) );
OR2XL U_g812 (.A(G2549_962_ngat), .B(G2546_743_ngat), .Y(G1551_1062_gat) );
AND5XL U_g813 (.A(G1584_993_gat), .B(G1588_990_gat), .C(G1592_987_gat), .D(G1596_984_gat), .E(G1600_981_gat), .Y(G1554_1063_gat) );
AND5XL U_g814 (.A(G1564_1008_gat), .B(G1568_1005_gat), .C(G1572_1002_gat), .D(G1576_999_gat), .E(G1580_996_gat), .Y(G1555_1064_gat) );
OR2XL U_g815 (.A(G2214_1025_ngat), .B(G2207_759_ngat), .Y(G2216_1065_gat) );
AND3XL U_g816 (.A(G1805_1016_gat), .B(G1767_925_gat), .C(G1754_854_gat), .Y(G1817_1066_gat) );
INVXL U_g817 (.A(G504_1012_gat), .Y(G505_1067_gat) );
INVXL U_g818 (.A(G731_1013_gat), .Y(G732_1068_gat) );
AND3XL U_g819 (.A(G1801_1017_gat), .B(G1763_857_gat), .C(G1758_924_gat), .Y(G1814_1069_gat) );
INVXL U_g820 (.A(G510_1014_gat), .Y(G511_1070_gat) );
INVXL U_g821 (.A(G737_1015_gat), .Y(G738_1071_gat) );
INVXL U_g822 (.A(G498_1019_gat), .Y(G499_1072_gat) );
INVXL U_g823 (.A(G725_1020_gat), .Y(G726_1073_gat) );
INVXL U_g824 (.A(G580_1023_gat), .Y(G584_1074_gat) );
BUFX20 U_g825 (.A(G610_1024_gat), .Y(G621_1075_gat) );
BUFX20 U_g826 (.A(G610_1024_gat), .Y(G625_1076_gat) );
BUFX20 U_g827 (.A(G589_1026_gat), .Y(G617_1077_gat) );
BUFX20 U_g828 (.A(G589_1026_gat), .Y(G613_1078_gat) );
INVXL U_g829 (.A(G2200_1031_gat), .Y(G2204_1079_gat) );
INVXL U_g830 (.A(G2220_1032_gat), .Y(G2224_1080_gat) );
INVXL U_g831 (.A(G2197_1033_gat), .Y(G2203_1081_gat) );
INVXL U_g832 (.A(G2217_1034_gat), .Y(G2223_1082_gat) );
INVXL U_g833 (.A(G492_1035_gat), .Y(G493_1083_gat) );
INVXL U_g834 (.A(G719_1036_gat), .Y(G720_1084_gat) );
AND2XL U_g835 (.A(G1845_953_gat), .B(G1874_975_gat), .Y(G1889_1085_gat) );
AND2XL U_g836 (.A(G1845_953_gat), .B(G1872_979_gat), .Y(G1887_1086_gat) );
AND2XL U_g837 (.A(G1845_953_gat), .B(G1870_982_gat), .Y(G1885_1087_gat) );
AND2XL U_g838 (.A(G1845_953_gat), .B(G1876_972_gat), .Y(G1891_1088_gat) );
AND2XL U_g839 (.A(G1907_954_gat), .B(G1936_976_gat), .Y(G1951_1089_gat) );
AND2XL U_g840 (.A(G1907_954_gat), .B(G1934_980_gat), .Y(G1949_1090_gat) );
AND2XL U_g841 (.A(G1907_954_gat), .B(G1932_983_gat), .Y(G1947_1091_gat) );
AND2XL U_g842 (.A(G1907_954_gat), .B(G1938_973_gat), .Y(G1953_1092_gat) );
AND2XL U_g843 (.A(G2062_968_gat), .B(G2065_715_gat), .Y(G1557_1093_gat) );
AND2XL U_g844 (.A(G1831_409_gat), .B(G1868_985_gat), .Y(G1883_1094_gat) );
AND2XL U_g845 (.A(G1831_409_gat), .B(G1866_988_gat), .Y(G1881_1095_gat) );
AND2XL U_g846 (.A(G1893_410_gat), .B(G1930_986_gat), .Y(G1945_1096_gat) );
AND2XL U_g847 (.A(G1893_410_gat), .B(G1928_989_gat), .Y(G1943_1097_gat) );
AND2XL U_g848 (.A(G748_411_gat), .B(G519_1027_gat), .Y(G521_1098_gat) );
AND2XL U_g849 (.A(G748_411_gat), .B(G525_1029_gat), .Y(G527_1099_gat) );
INVXL U_g850 (.A(G533_1041_gat), .Y(G534_1100_gat) );
INVXL U_g851 (.A(G539_1042_gat), .Y(G540_1101_gat) );
AND2XL U_g852 (.A(G994_412_gat), .B(G693_1028_gat), .Y(G695_1102_gat) );
AND2XL U_g853 (.A(G994_412_gat), .B(G699_1030_gat), .Y(G701_1103_gat) );
INVXL U_g854 (.A(G707_1043_gat), .Y(G708_1104_gat) );
INVXL U_g855 (.A(G713_1044_gat), .Y(G714_1105_gat) );
INVXL U_g856 (.A(G1091_1045_gat), .Y(G1092_1106_gat) );
INVXL U_g857 (.A(G2722_1047_gat), .Y(G2726_1107_gat) );
OR2XL U_g858 (.A(G1829_966_ngat), .B(G1828_1048_ngat), .Y(G1830_1108_gat) );
AND2XL U_g859 (.A(G1558_1053_gat), .B(G1557_1093_gat), .Y(G1559_1109_gat) );
OR2XL U_g860 (.A(G1552_978_ngat), .B(G1551_1062_ngat), .Y(G1553_1110_gat) );
AND2XL U_g861 (.A(G1555_1064_gat), .B(G1554_1063_gat), .Y(G1556_1111_gat) );
OR2XL U_g862 (.A(G1863_991_gat), .B(G1861_1049_gat), .Y(G1864_1112_gat) );
OR2XL U_g863 (.A(G1925_992_gat), .B(G1923_1050_gat), .Y(G1926_1113_gat) );
OR2XL U_g864 (.A(G1858_994_gat), .B(G1856_1051_gat), .Y(G1859_1114_gat) );
OR2XL U_g865 (.A(G1920_995_gat), .B(G1918_1052_gat), .Y(G1921_1115_gat) );
OR2XL U_g866 (.A(G1377_997_gat), .B(G1375_1054_gat), .Y(G1382_1116_gat) );
OR2XL U_g867 (.A(G1623_998_gat), .B(G1621_1055_gat), .Y(G1628_1117_gat) );
OR2XL U_g868 (.A(G1373_1000_gat), .B(G1371_1056_gat), .Y(G1380_1118_gat) );
OR2XL U_g869 (.A(G1619_1001_gat), .B(G1617_1057_gat), .Y(G1626_1119_gat) );
OR2XL U_g870 (.A(G1615_1003_gat), .B(G1614_1059_gat), .Y(G1624_1120_gat) );
OR2XL U_g871 (.A(G1369_1004_gat), .B(G1368_1058_gat), .Y(G1378_1121_gat) );
OR2XL U_g872 (.A(G676_1006_gat), .B(G675_1060_gat), .Y(G677_1122_gat) );
OR2XL U_g873 (.A(G1108_1007_gat), .B(G1107_1061_gat), .Y(G1109_1123_gat) );
OR2XL U_g874 (.A(G2216_1065_ngat), .B(G2215_1009_ngat), .Y(G2238_1124_gat) );
AND3XL U_g875 (.A(G621_1075_gat), .B(G592_760_gat), .C(G601_930_gat), .Y(G636_1125_gat) );
AND3XL U_g876 (.A(G625_1076_gat), .B(G596_853_gat), .C(G605_1022_gat), .Y(G639_1126_gat) );
AND2XL U_g877 (.A(G1815_1010_ngat), .B(G1814_1069_ngat), .Y(G1816_1127_gat) );
AND2XL U_g878 (.A(G1818_1011_ngat), .B(G1817_1066_ngat), .Y(G1819_1128_gat) );
AND2XL U_g879 (.A(G505_1067_gat), .B(G1889_1085_gat), .Y(G915_1129_gat) );
BUFX20 U_g880 (.A(G505_1067_gat), .Y(G2278_1130_gat) );
AND2XL U_g881 (.A(G732_1068_gat), .B(G1951_1089_gat), .Y(G1133_1131_gat) );
BUFX20 U_g882 (.A(G732_1068_gat), .Y(G2366_1132_gat) );
AND2XL U_g883 (.A(G511_1070_gat), .B(G1891_1088_gat), .Y(G907_1133_gat) );
BUFX20 U_g884 (.A(G511_1070_gat), .Y(G2270_1134_gat) );
AND2XL U_g885 (.A(G738_1071_gat), .B(G1953_1092_gat), .Y(G1125_1135_gat) );
BUFX20 U_g886 (.A(G738_1071_gat), .Y(G2358_1136_gat) );
AND2XL U_g887 (.A(G499_1072_gat), .B(G1887_1086_gat), .Y(G922_1137_gat) );
BUFX20 U_g888 (.A(G499_1072_gat), .Y(G2286_1138_gat) );
AND2XL U_g889 (.A(G726_1073_gat), .B(G1949_1090_gat), .Y(G1140_1139_gat) );
BUFX20 U_g890 (.A(G726_1073_gat), .Y(G2374_1140_gat) );
AND3XL U_g891 (.A(G613_1078_gat), .B(G571_929_gat), .C(G580_1023_gat), .Y(G630_1141_gat) );
AND3XL U_g892 (.A(G617_1077_gat), .B(G575_1021_gat), .C(G584_1074_gat), .Y(G633_1142_gat) );
INVXL U_g893 (.A(G621_1075_gat), .Y(G624_1143_gat) );
INVXL U_g894 (.A(G625_1076_gat), .Y(G628_1144_gat) );
INVXL U_g895 (.A(G617_1077_gat), .Y(G620_1145_gat) );
INVXL U_g896 (.A(G613_1078_gat), .Y(G616_1146_gat) );
OR2XL U_g897 (.A(G2203_1081_ngat), .B(G2200_1031_ngat), .Y(G2205_1147_gat) );
OR2XL U_g898 (.A(G2223_1082_ngat), .B(G2220_1032_ngat), .Y(G2225_1148_gat) );
OR2XL U_g899 (.A(G2204_1079_ngat), .B(G2197_1033_ngat), .Y(G2206_1149_gat) );
OR2XL U_g900 (.A(G2224_1080_ngat), .B(G2217_1034_ngat), .Y(G2226_1150_gat) );
AND2XL U_g901 (.A(G1885_1087_gat), .B(G493_1083_gat), .Y(G924_1151_gat) );
BUFX20 U_g902 (.A(G493_1083_gat), .Y(G2294_1152_gat) );
AND2XL U_g903 (.A(G1947_1091_gat), .B(G720_1084_gat), .Y(G1142_1153_gat) );
BUFX20 U_g904 (.A(G720_1084_gat), .Y(G2382_1154_gat) );
BUFX20 U_g905 (.A(G1889_1085_gat), .Y(G2275_1155_gat) );
BUFX20 U_g906 (.A(G1887_1086_gat), .Y(G2283_1156_gat) );
BUFX20 U_g907 (.A(G1885_1087_gat), .Y(G2291_1157_gat) );
BUFX20 U_g908 (.A(G1891_1088_gat), .Y(G2267_1158_gat) );
BUFX20 U_g909 (.A(G1951_1089_gat), .Y(G2363_1159_gat) );
BUFX20 U_g910 (.A(G1949_1090_gat), .Y(G2371_1160_gat) );
BUFX20 U_g911 (.A(G1947_1091_gat), .Y(G2379_1161_gat) );
BUFX20 U_g912 (.A(G1953_1092_gat), .Y(G2355_1162_gat) );
AND2XL U_g913 (.A(G540_1101_gat), .B(G1883_1094_gat), .Y(G937_1163_gat) );
BUFX20 U_g914 (.A(G1883_1094_gat), .Y(G2299_1164_gat) );
AND2XL U_g915 (.A(G534_1100_gat), .B(G1881_1095_gat), .Y(G946_1165_gat) );
BUFX20 U_g916 (.A(G1881_1095_gat), .Y(G2307_1166_gat) );
AND2XL U_g917 (.A(G714_1105_gat), .B(G1945_1096_gat), .Y(G1155_1167_gat) );
BUFX20 U_g918 (.A(G1945_1096_gat), .Y(G2387_1168_gat) );
AND2XL U_g919 (.A(G708_1104_gat), .B(G1943_1097_gat), .Y(G1164_1169_gat) );
BUFX20 U_g920 (.A(G1943_1097_gat), .Y(G2395_1170_gat) );
INVXL U_g921 (.A(G521_1098_gat), .Y(G522_1171_gat) );
INVXL U_g922 (.A(G527_1099_gat), .Y(G528_1172_gat) );
BUFX20 U_g923 (.A(G534_1100_gat), .Y(G2310_1173_gat) );
BUFX20 U_g924 (.A(G540_1101_gat), .Y(G2302_1174_gat) );
INVXL U_g925 (.A(G695_1102_gat), .Y(G696_1175_gat) );
INVXL U_g926 (.A(G701_1103_gat), .Y(G702_1176_gat) );
BUFX20 U_g927 (.A(G708_1104_gat), .Y(G2398_1177_gat) );
BUFX20 U_g928 (.A(G714_1105_gat), .Y(G2390_1178_gat) );
BUFX20 U_g929 (.A(G1382_1116_gat), .Y(G2331_1181_gat) );
BUFX20 U_g930 (.A(G1628_1117_gat), .Y(G2419_1182_gat) );
BUFX20 U_g931 (.A(G1380_1118_gat), .Y(G2251_1183_gat) );
BUFX20 U_g932 (.A(G1626_1119_gat), .Y(G2339_1184_gat) );
BUFX20 U_g933 (.A(G1624_1120_gat), .Y(G2347_1185_gat) );
BUFX20 U_g934 (.A(G1378_1121_gat), .Y(G2259_1186_gat) );
INVXL U_g935 (.A(G2238_1124_gat), .Y(G2242_1187_gat) );
AND3XL U_g936 (.A(G628_1144_gat), .B(G605_1022_gat), .C(G592_760_gat), .Y(G638_1188_gat) );
AND3XL U_g937 (.A(G624_1143_gat), .B(G601_930_gat), .C(G596_853_gat), .Y(G635_1189_gat) );
OR2XL U_g938 (.A(G1816_1127_ngat), .B(G1819_1128_ngat), .Y(G2719_1190_gat) );
INVXL U_g939 (.A(G2278_1130_gat), .Y(G2282_1191_gat) );
INVXL U_g940 (.A(G2366_1132_gat), .Y(G2370_1192_gat) );
INVXL U_g941 (.A(G2270_1134_gat), .Y(G2274_1193_gat) );
INVXL U_g942 (.A(G2358_1136_gat), .Y(G2362_1194_gat) );
INVXL U_g943 (.A(G2286_1138_gat), .Y(G2290_1195_gat) );
INVXL U_g944 (.A(G2374_1140_gat), .Y(G2378_1196_gat) );
OR2XL U_g945 (.A(G2241_770_ngat), .B(G2238_1124_ngat), .Y(G645_1197_gat) );
AND3XL U_g946 (.A(G620_1145_gat), .B(G584_1074_gat), .C(G571_929_gat), .Y(G632_1198_gat) );
AND3XL U_g947 (.A(G616_1146_gat), .B(G580_1023_gat), .C(G575_1021_gat), .Y(G629_1199_gat) );
AND2XL U_g948 (.A(G1035_618_gat), .B(G1378_1121_gat), .Y(G674_1200_gat) );
AND2XL U_g949 (.A(G1035_618_gat), .B(G1624_1120_gat), .Y(G1106_1201_gat) );
AND2XL U_g950 (.A(G1043_693_gat), .B(G1380_1118_gat), .Y(G671_1202_gat) );
AND2XL U_g951 (.A(G1043_693_gat), .B(G1626_1119_gat), .Y(G1104_1203_gat) );
AND2XL U_g952 (.A(G1051_695_gat), .B(G1382_1116_gat), .Y(G967_1204_gat) );
AND2XL U_g953 (.A(G1051_695_gat), .B(G1628_1117_gat), .Y(G1184_1205_gat) );
OR2XL U_g954 (.A(G2206_1149_ngat), .B(G2205_1147_ngat), .Y(G2230_1206_gat) );
OR2XL U_g955 (.A(G2226_1150_ngat), .B(G2225_1148_ngat), .Y(G2246_1207_gat) );
INVXL U_g956 (.A(G2294_1152_gat), .Y(G2298_1208_gat) );
INVXL U_g957 (.A(G2382_1154_gat), .Y(G2386_1209_gat) );
AND2XL U_g958 (.A(G1031_630_gat), .B(G677_1122_gat), .Y(G679_1210_gat) );
AND2XL U_g959 (.A(G1031_630_gat), .B(G1109_1123_gat), .Y(G1110_1211_gat) );
INVXL U_g960 (.A(G2275_1155_gat), .Y(G2281_1212_gat) );
INVXL U_g961 (.A(G2283_1156_gat), .Y(G2289_1213_gat) );
INVXL U_g962 (.A(G2291_1157_gat), .Y(G2297_1214_gat) );
INVXL U_g963 (.A(G2267_1158_gat), .Y(G2273_1215_gat) );
INVXL U_g964 (.A(G2363_1159_gat), .Y(G2369_1216_gat) );
INVXL U_g965 (.A(G2371_1160_gat), .Y(G2377_1217_gat) );
INVXL U_g966 (.A(G2379_1161_gat), .Y(G2385_1218_gat) );
INVXL U_g967 (.A(G2355_1162_gat), .Y(G2361_1219_gat) );
AND2XL U_g968 (.A(G14_9_gat), .B(G1092_1106_gat), .Y(G401_1276_gat) );
AND3XL U_g969 (.A(G894_533_gat), .B(G1559_1109_gat), .C(G1556_1111_gat), .Y(G311_1278_gat) );
INVXL U_g970 (.A(G2299_1164_gat), .Y(G2305_1222_gat) );
INVXL U_g971 (.A(G2307_1166_gat), .Y(G2313_1223_gat) );
AND2XL U_g972 (.A(G1831_409_gat), .B(G1864_1112_gat), .Y(G1879_1224_gat) );
AND2XL U_g973 (.A(G1831_409_gat), .B(G1859_1114_gat), .Y(G1877_1225_gat) );
INVXL U_g974 (.A(G2387_1168_gat), .Y(G2393_1226_gat) );
INVXL U_g975 (.A(G2395_1170_gat), .Y(G2401_1227_gat) );
AND2XL U_g976 (.A(G1893_410_gat), .B(G1926_1113_gat), .Y(G1941_1228_gat) );
AND2XL U_g977 (.A(G1893_410_gat), .B(G1921_1115_gat), .Y(G1939_1229_gat) );
BUFX20 U_g978 (.A(G522_1171_gat), .Y(G2326_1230_gat) );
BUFX20 U_g979 (.A(G528_1172_gat), .Y(G2318_1231_gat) );
INVXL U_g980 (.A(G2310_1173_gat), .Y(G2314_1232_gat) );
INVXL U_g981 (.A(G2302_1174_gat), .Y(G2306_1233_gat) );
BUFX20 U_g982 (.A(G696_1175_gat), .Y(G2414_1234_gat) );
BUFX20 U_g983 (.A(G702_1176_gat), .Y(G2406_1235_gat) );
INVXL U_g984 (.A(G2398_1177_gat), .Y(G2402_1236_gat) );
INVXL U_g985 (.A(G2390_1178_gat), .Y(G2394_1237_gat) );
OR2XL U_g986 (.A(G2726_1107_ngat), .B(G2719_1190_ngat), .Y(G1827_1238_gat) );
INVXL U_g987 (.A(G2331_1181_gat), .Y(G2337_1239_gat) );
INVXL U_g988 (.A(G2419_1182_gat), .Y(G2425_1240_gat) );
INVXL U_g989 (.A(G2251_1183_gat), .Y(G2257_1241_gat) );
INVXL U_g990 (.A(G2339_1184_gat), .Y(G2345_1242_gat) );
INVXL U_g991 (.A(G2347_1185_gat), .Y(G2353_1243_gat) );
INVXL U_g992 (.A(G2259_1186_gat), .Y(G2265_1244_gat) );
AND2XL U_g993 (.A(G636_1125_ngat), .B(G635_1189_ngat), .Y(G637_1245_gat) );
AND2XL U_g994 (.A(G639_1126_ngat), .B(G638_1188_ngat), .Y(G640_1246_gat) );
INVXL U_g995 (.A(G2719_1190_gat), .Y(G2725_1247_gat) );
OR2XL U_g996 (.A(G2281_1212_ngat), .B(G2278_1130_ngat), .Y(G908_1248_gat) );
OR2XL U_g997 (.A(G2369_1216_ngat), .B(G2366_1132_ngat), .Y(G1126_1249_gat) );
OR2XL U_g998 (.A(G2273_1215_ngat), .B(G2270_1134_ngat), .Y(G899_1250_gat) );
OR2XL U_g999 (.A(G2361_1219_ngat), .B(G2358_1136_ngat), .Y(G1117_1251_gat) );
OR2XL U_g1000 (.A(G2289_1213_ngat), .B(G2286_1138_ngat), .Y(G916_1252_gat) );
OR2XL U_g1001 (.A(G2377_1217_ngat), .B(G2374_1140_ngat), .Y(G1134_1253_gat) );
OR2XL U_g1002 (.A(G2242_1187_ngat), .B(G2235_684_ngat), .Y(G646_1254_gat) );
AND2XL U_g1003 (.A(G630_1141_ngat), .B(G629_1199_ngat), .Y(G631_1255_gat) );
AND2XL U_g1004 (.A(G633_1142_ngat), .B(G632_1198_ngat), .Y(G634_1256_gat) );
OR2XL U_g1005 (.A(G2354_773_ngat), .B(G2347_1185_ngat), .Y(G1115_1257_gat) );
OR2XL U_g1006 (.A(G2266_775_ngat), .B(G2259_1186_ngat), .Y(G684_1258_gat) );
OR2XL U_g1007 (.A(G2346_868_ngat), .B(G2339_1184_ngat), .Y(G1099_1259_gat) );
OR2XL U_g1008 (.A(G2258_870_ngat), .B(G2251_1183_ngat), .Y(G665_1260_gat) );
OR2XL U_g1009 (.A(G2426_872_ngat), .B(G2419_1182_ngat), .Y(G1181_1261_gat) );
OR2XL U_g1010 (.A(G2338_873_ngat), .B(G2331_1181_ngat), .Y(G963_1262_gat) );
INVXL U_g1011 (.A(G2230_1206_gat), .Y(G2234_1263_gat) );
INVXL U_g1012 (.A(G2246_1207_gat), .Y(G2250_1264_gat) );
OR2XL U_g1013 (.A(G2297_1214_ngat), .B(G2294_1152_ngat), .Y(G925_1265_gat) );
OR2XL U_g1014 (.A(G2385_1218_ngat), .B(G2382_1154_ngat), .Y(G1143_1266_gat) );
OR2XL U_g1015 (.A(G2282_1191_ngat), .B(G2275_1155_ngat), .Y(G909_1267_gat) );
OR2XL U_g1016 (.A(G2290_1195_ngat), .B(G2283_1156_ngat), .Y(G917_1268_gat) );
OR2XL U_g1017 (.A(G2298_1208_ngat), .B(G2291_1157_ngat), .Y(G926_1269_gat) );
OR2XL U_g1018 (.A(G2274_1193_ngat), .B(G2267_1158_ngat), .Y(G900_1270_gat) );
OR2XL U_g1019 (.A(G2370_1192_ngat), .B(G2363_1159_ngat), .Y(G1127_1271_gat) );
OR2XL U_g1020 (.A(G2378_1196_ngat), .B(G2371_1160_ngat), .Y(G1135_1272_gat) );
OR2XL U_g1021 (.A(G2386_1209_ngat), .B(G2379_1161_ngat), .Y(G1144_1273_gat) );
OR2XL U_g1022 (.A(G2362_1194_ngat), .B(G2355_1162_ngat), .Y(G1118_1274_gat) );
INVXL U_g1023 (.A(G401_1276_gat), .Y(G1087_1275_gat) );
OR2XL U_g1024 (.A(G2306_1233_ngat), .B(G2299_1164_ngat), .Y(G929_1279_gat) );
OR2XL U_g1025 (.A(G2314_1232_ngat), .B(G2307_1166_ngat), .Y(G939_1280_gat) );
BUFX20 U_g1026 (.A(G1879_1224_gat), .Y(G2315_1281_gat) );
BUFX20 U_g1027 (.A(G1877_1225_gat), .Y(G2323_1282_gat) );
OR2XL U_g1028 (.A(G2394_1237_ngat), .B(G2387_1168_ngat), .Y(G1147_1283_gat) );
OR2XL U_g1029 (.A(G2402_1236_ngat), .B(G2395_1170_ngat), .Y(G1157_1284_gat) );
BUFX20 U_g1030 (.A(G1941_1228_gat), .Y(G2403_1285_gat) );
BUFX20 U_g1031 (.A(G1939_1229_gat), .Y(G2411_1286_gat) );
INVXL U_g1032 (.A(G2326_1230_gat), .Y(G2330_1287_gat) );
AND2XL U_g1033 (.A(G522_1171_gat), .B(G1877_1225_gat), .Y(G961_1288_gat) );
AND2XL U_g1034 (.A(G528_1172_gat), .B(G1879_1224_gat), .Y(G954_1289_gat) );
INVXL U_g1035 (.A(G2318_1231_gat), .Y(G2322_1290_gat) );
OR2XL U_g1036 (.A(G2313_1223_ngat), .B(G2310_1173_ngat), .Y(G938_1291_gat) );
OR2XL U_g1037 (.A(G2305_1222_ngat), .B(G2302_1174_ngat), .Y(G928_1292_gat) );
INVXL U_g1038 (.A(G2414_1234_gat), .Y(G2418_1293_gat) );
AND2XL U_g1039 (.A(G696_1175_gat), .B(G1939_1229_gat), .Y(G1179_1294_gat) );
AND2XL U_g1040 (.A(G702_1176_gat), .B(G1941_1228_gat), .Y(G1172_1295_gat) );
INVXL U_g1041 (.A(G2406_1235_gat), .Y(G2410_1296_gat) );
OR2XL U_g1042 (.A(G2401_1227_ngat), .B(G2398_1177_ngat), .Y(G1156_1297_gat) );
OR2XL U_g1043 (.A(G2393_1226_ngat), .B(G2390_1178_ngat), .Y(G1146_1298_gat) );
OR2XL U_g1044 (.A(G2725_1247_ngat), .B(G2722_1047_ngat), .Y(G1826_1299_gat) );
OR2XL U_g1045 (.A(G637_1245_ngat), .B(G640_1246_ngat), .Y(G2243_1300_gat) );
OR2XL U_g1046 (.A(G909_1267_ngat), .B(G908_1248_ngat), .Y(G910_1301_gat) );
OR2XL U_g1047 (.A(G1127_1271_ngat), .B(G1126_1249_ngat), .Y(G1128_1302_gat) );
OR2XL U_g1048 (.A(G900_1270_ngat), .B(G899_1250_ngat), .Y(G901_1303_gat) );
OR2XL U_g1049 (.A(G1118_1274_ngat), .B(G1117_1251_ngat), .Y(G1119_1304_gat) );
OR2XL U_g1050 (.A(G917_1268_ngat), .B(G916_1252_ngat), .Y(G918_1305_gat) );
OR2XL U_g1051 (.A(G1135_1272_ngat), .B(G1134_1253_ngat), .Y(G1136_1306_gat) );
OR2XL U_g1052 (.A(G646_1254_ngat), .B(G645_1197_ngat), .Y(G647_1307_gat) );
OR2XL U_g1053 (.A(G631_1255_ngat), .B(G634_1256_ngat), .Y(G2227_1308_gat) );
OR2XL U_g1054 (.A(G2353_1243_ngat), .B(G2350_687_ngat), .Y(G1114_1309_gat) );
OR2XL U_g1055 (.A(G2265_1244_ngat), .B(G2262_689_ngat), .Y(G683_1310_gat) );
OR2XL U_g1056 (.A(G2345_1242_ngat), .B(G2342_779_ngat), .Y(G1098_1311_gat) );
OR2XL U_g1057 (.A(G2257_1241_ngat), .B(G2254_781_ngat), .Y(G664_1312_gat) );
OR2XL U_g1058 (.A(G2425_1240_ngat), .B(G2422_783_ngat), .Y(G1180_1313_gat) );
OR2XL U_g1059 (.A(G2337_1239_ngat), .B(G2334_784_ngat), .Y(G962_1314_gat) );
OR2XL U_g1060 (.A(G926_1269_ngat), .B(G925_1265_ngat), .Y(G927_1315_gat) );
OR2XL U_g1061 (.A(G1144_1273_ngat), .B(G1143_1266_ngat), .Y(G1145_1316_gat) );
OR2XL U_g1062 (.A(G929_1279_ngat), .B(G928_1292_ngat), .Y(G930_1317_gat) );
OR2XL U_g1063 (.A(G939_1280_ngat), .B(G938_1291_ngat), .Y(G940_1318_gat) );
OR2XL U_g1064 (.A(G2322_1290_ngat), .B(G2315_1281_ngat), .Y(G948_1319_gat) );
INVXL U_g1065 (.A(G2315_1281_gat), .Y(G2321_1320_gat) );
OR2XL U_g1066 (.A(G2330_1287_ngat), .B(G2323_1282_ngat), .Y(G956_1321_gat) );
INVXL U_g1067 (.A(G2323_1282_gat), .Y(G2329_1322_gat) );
OR2XL U_g1068 (.A(G1147_1283_ngat), .B(G1146_1298_ngat), .Y(G1148_1323_gat) );
OR2XL U_g1069 (.A(G1157_1284_ngat), .B(G1156_1297_ngat), .Y(G1158_1324_gat) );
OR2XL U_g1070 (.A(G2410_1296_ngat), .B(G2403_1285_ngat), .Y(G1166_1325_gat) );
INVXL U_g1071 (.A(G2403_1285_gat), .Y(G2409_1326_gat) );
OR2XL U_g1072 (.A(G2418_1293_ngat), .B(G2411_1286_ngat), .Y(G1174_1327_gat) );
INVXL U_g1073 (.A(G2411_1286_gat), .Y(G2417_1328_gat) );
OR2XL U_g1074 (.A(G1827_1238_ngat), .B(G1826_1299_ngat), .Y(G686_1329_gat) );
AND2XL U_g1075 (.A(G865_291_gat), .B(G647_1307_gat), .Y(G143_1330_gat) );
INVXL U_g1076 (.A(G2243_1300_gat), .Y(G2249_1331_gat) );
AND2XL U_g1077 (.A(G915_1129_gat), .B(G901_1303_gat), .Y(G970_1332_gat) );
AND4XL U_g1078 (.A(G901_1303_gat), .B(G918_1305_gat), .C(G927_1315_gat), .D(G910_1301_gat), .Y(G968_1333_gat) );
AND2XL U_g1079 (.A(G1133_1131_gat), .B(G1119_1304_gat), .Y(G1187_1334_gat) );
AND4XL U_g1080 (.A(G1119_1304_gat), .B(G1136_1306_gat), .C(G1145_1316_gat), .D(G1128_1302_gat), .Y(G1185_1335_gat) );
AND3XL U_g1081 (.A(G922_1137_gat), .B(G901_1303_gat), .C(G910_1301_gat), .Y(G971_1336_gat) );
AND3XL U_g1082 (.A(G1140_1139_gat), .B(G1119_1304_gat), .C(G1128_1302_gat), .Y(G1188_1337_gat) );
INVXL U_g1083 (.A(G2227_1308_gat), .Y(G2233_1338_gat) );
OR2XL U_g1084 (.A(G1115_1257_ngat), .B(G1114_1309_ngat), .Y(G1112_1339_gat) );
OR2XL U_g1085 (.A(G684_1258_ngat), .B(G683_1310_ngat), .Y(G681_1340_gat) );
OR2XL U_g1086 (.A(G1099_1259_ngat), .B(G1098_1311_ngat), .Y(G1100_1341_gat) );
OR2XL U_g1087 (.A(G665_1260_ngat), .B(G664_1312_ngat), .Y(G666_1342_gat) );
OR2XL U_g1088 (.A(G1181_1261_ngat), .B(G1180_1313_ngat), .Y(G1182_1343_gat) );
OR2XL U_g1089 (.A(G963_1262_ngat), .B(G962_1314_ngat), .Y(G964_1344_gat) );
OR2XL U_g1090 (.A(G2234_1263_ngat), .B(G2227_1308_ngat), .Y(G642_1345_gat) );
OR2XL U_g1091 (.A(G2250_1264_ngat), .B(G2243_1300_ngat), .Y(G649_1346_gat) );
AND4XL U_g1092 (.A(G910_1301_gat), .B(G924_1151_gat), .C(G901_1303_gat), .D(G918_1305_gat), .Y(G972_1347_gat) );
AND4XL U_g1093 (.A(G1128_1302_gat), .B(G1142_1153_gat), .C(G1119_1304_gat), .D(G1136_1306_gat), .Y(G1189_1348_gat) );
AND2XL U_g1094 (.A(G946_1165_gat), .B(G930_1317_gat), .Y(G978_1349_gat) );
AND2XL U_g1095 (.A(G1164_1169_gat), .B(G1148_1323_gat), .Y(G1195_1350_gat) );
OR2XL U_g1096 (.A(G2329_1322_ngat), .B(G2326_1230_ngat), .Y(G955_1351_gat) );
AND3XL U_g1097 (.A(G954_1289_gat), .B(G930_1317_gat), .C(G940_1318_gat), .Y(G979_1352_gat) );
OR2XL U_g1098 (.A(G2321_1320_ngat), .B(G2318_1231_ngat), .Y(G947_1353_gat) );
OR2XL U_g1099 (.A(G2417_1328_ngat), .B(G2414_1234_ngat), .Y(G1173_1354_gat) );
AND3XL U_g1100 (.A(G1172_1295_gat), .B(G1148_1323_gat), .C(G1158_1324_gat), .Y(G1196_1355_gat) );
OR2XL U_g1101 (.A(G2409_1326_ngat), .B(G2406_1235_ngat), .Y(G1165_1356_gat) );
INVXL U_g1102 (.A(G686_1329_gat), .Y(G687_1357_gat) );
INVXL U_g1103 (.A(G968_1333_gat), .Y(G969_1359_gat) );
INVXL U_g1104 (.A(G1185_1335_gat), .Y(G1186_1360_gat) );
OR4XL U_g1105 (.A(G972_1347_gat), .B(G971_1336_gat), .C(G970_1332_gat), .D(G907_1133_gat), .Y(G973_1361_gat) );
OR4XL U_g1106 (.A(G1189_1348_gat), .B(G1188_1337_gat), .C(G1187_1334_gat), .D(G1125_1135_gat), .Y(G1190_1362_gat) );
AND2XL U_g1107 (.A(G674_1200_gat), .B(G666_1342_gat), .Y(G680_1363_gat) );
AND2XL U_g1108 (.A(G1106_1201_gat), .B(G1100_1341_gat), .Y(G1111_1364_gat) );
OR2XL U_g1109 (.A(G2233_1338_ngat), .B(G2230_1206_ngat), .Y(G641_1365_gat) );
OR2XL U_g1110 (.A(G2249_1331_ngat), .B(G2246_1207_ngat), .Y(G648_1366_gat) );
AND3XL U_g1111 (.A(G679_1210_gat), .B(G666_1342_gat), .C(G681_1340_gat), .Y(G682_1367_gat) );
AND3XL U_g1112 (.A(G1110_1211_gat), .B(G1100_1341_gat), .C(G1112_1339_gat), .Y(G1113_1368_gat) );
OR2XL U_g1113 (.A(G948_1319_ngat), .B(G947_1353_ngat), .Y(G949_1369_gat) );
OR2XL U_g1114 (.A(G956_1321_ngat), .B(G955_1351_ngat), .Y(G957_1370_gat) );
OR2XL U_g1115 (.A(G1166_1325_ngat), .B(G1165_1356_ngat), .Y(G1167_1371_gat) );
OR2XL U_g1116 (.A(G1174_1327_ngat), .B(G1173_1354_ngat), .Y(G1175_1372_gat) );
INVXL U_g1117 (.A(G973_1361_gat), .Y(G976_1373_gat) );
INVXL U_g1118 (.A(G1190_1362_gat), .Y(G1193_1374_gat) );
OR3XL U_g1119 (.A(G682_1367_gat), .B(G680_1363_gat), .C(G671_1202_gat), .Y(G685_1375_gat) );
OR3XL U_g1120 (.A(G1113_1368_gat), .B(G1111_1364_gat), .C(G1104_1203_gat), .Y(G1116_1376_gat) );
AND5XL U_g1121 (.A(G940_1318_gat), .B(G967_1204_gat), .C(G930_1317_gat), .D(G949_1369_gat), .E(G957_1370_gat), .Y(G981_1377_gat) );
AND5XL U_g1122 (.A(G1158_1324_gat), .B(G1184_1205_gat), .C(G1148_1323_gat), .D(G1167_1371_gat), .E(G1175_1372_gat), .Y(G1198_1378_gat) );
OR2XL U_g1123 (.A(G642_1345_ngat), .B(G641_1365_ngat), .Y(G643_1379_gat) );
OR2XL U_g1124 (.A(G649_1346_ngat), .B(G648_1366_ngat), .Y(G650_1380_gat) );
AND2XL U_g1125 (.A(G487_403_gat), .B(G687_1357_gat), .Y(G395_1392_gat) );
AND5XL U_g1126 (.A(G957_1370_gat), .B(G930_1317_gat), .C(G949_1369_gat), .D(G964_1344_gat), .E(G940_1318_gat), .Y(G977_1382_gat) );
AND5XL U_g1127 (.A(G1175_1372_gat), .B(G1148_1323_gat), .C(G1167_1371_gat), .D(G1182_1343_gat), .E(G1158_1324_gat), .Y(G1194_1383_gat) );
AND4XL U_g1128 (.A(G940_1318_gat), .B(G961_1288_gat), .C(G930_1317_gat), .D(G949_1369_gat), .Y(G980_1384_gat) );
AND4XL U_g1129 (.A(G1158_1324_gat), .B(G1179_1294_gat), .C(G1148_1323_gat), .D(G1167_1371_gat), .Y(G1197_1385_gat) );
AND2XL U_g1130 (.A(G868_198_gat), .B(G650_1380_gat), .Y(G884_1386_gat) );
OR2XL U_g1131 (.A(G969_1359_ngat), .B(G976_1373_ngat), .Y(G988_1387_gat) );
OR2XL U_g1132 (.A(G1186_1360_ngat), .B(G1193_1374_ngat), .Y(G1205_1388_gat) );
AND2XL U_g1133 (.A(G685_1375_gat), .B(G977_1382_gat), .Y(G983_1389_gat) );
AND2XL U_g1134 (.A(G1116_1376_gat), .B(G1194_1383_gat), .Y(G1200_1390_gat) );
INVXL U_g1135 (.A(G643_1379_gat), .Y(G644_1391_gat) );
INVXL U_g1136 (.A(G395_1392_gat), .Y(G690_1393_gat) );
OR5XL U_g1137 (.A(G981_1377_gat), .B(G980_1384_gat), .C(G979_1352_gat), .D(G978_1349_gat), .E(G937_1163_gat), .Y(G982_1394_gat) );
OR5XL U_g1138 (.A(G1198_1378_gat), .B(G1197_1385_gat), .C(G1196_1355_gat), .D(G1195_1350_gat), .E(G1155_1167_gat), .Y(G1199_1395_gat) );
OR2XL U_g1139 (.A(G884_1386_gat), .B(G883_668_gat), .Y(G895_1396_gat) );
OR2XL U_g1140 (.A(G983_1389_gat), .B(G982_1394_gat), .Y(G984_1397_gat) );
OR2XL U_g1141 (.A(G1200_1390_gat), .B(G1199_1395_gat), .Y(G1201_1398_gat) );
AND2XL U_g1142 (.A(G487_403_gat), .B(G644_1391_gat), .Y(G397_1406_gat) );
AND2XL U_g1143 (.A(G984_1397_gat), .B(G988_1387_gat), .Y(G990_1402_gat) );
AND2XL U_g1144 (.A(G1201_1398_gat), .B(G1205_1388_gat), .Y(G1207_1403_gat) );
INVXL U_g1145 (.A(G984_1397_gat), .Y(G987_1404_gat) );
INVXL U_g1146 (.A(G1201_1398_gat), .Y(G1204_1405_gat) );
INVXL U_g1147 (.A(G397_1406_gat), .Y(G1027_1407_gat) );
AND3XL U_g1148 (.A(G1830_1108_gat), .B(G1027_1407_gat), .C(G690_1393_gat), .Y(G1085_1408_gat) );
AND2XL U_g1149 (.A(G987_1404_gat), .B(G973_1361_gat), .Y(G989_1409_gat) );
AND2XL U_g1150 (.A(G1204_1405_gat), .B(G1190_1362_gat), .Y(G1206_1410_gat) );
OR2XL U_g1151 (.A(G990_1402_gat), .B(G989_1409_gat), .Y(G991_1411_gat) );
OR2XL U_g1152 (.A(G1207_1403_gat), .B(G1206_1410_gat), .Y(G329_1414_gat) );
OR2XL U_g1153 (.A(G991_1411_ngat), .B(G329_1414_ngat), .Y(G1221_1413_gat) );
AND2XL U_g1154 (.A(G991_1411_gat), .B(G1221_1413_gat), .Y(G1239_1415_gat) );
AND2XL U_g1155 (.A(G1221_1413_gat), .B(G329_1414_gat), .Y(G1238_1416_gat) );
OR2XL U_g1156 (.A(G1239_1415_gat), .B(G1238_1416_gat), .Y(G1240_1417_gat) );
INVXL U_g1157 (.A(G1240_1417_gat), .Y(G1247_1418_gat) );
AND2XL U_g1158 (.A(G1247_1418_gat), .B(G1240_1417_gat), .Y(G471_1419_gat) );
OR2XL U_g1159 (.A(G1247_1418_gat), .B(G471_1419_gat), .Y(G473_1420_gat) );
AND3XL U_g1160 (.A(G473_1420_gat), .B(G1087_1275_gat), .C(G1553_1110_gat), .Y(G1088_1421_gat) );
AND3XL U_g1161 (.A(G319_656_gat), .B(G1088_1421_gat), .C(G1085_1408_gat), .Y(G308_1425_gat) );
BUFX20 U_g1162 (.A(GIN_169_114_gat), .Y(G169_114_gat) );
BUFX20 U_g1163 (.A(GIN_174_115_gat), .Y(G174_115_gat) );
BUFX20 U_g1164 (.A(GIN_177_116_gat), .Y(G177_116_gat) );
BUFX20 U_g1165 (.A(GIN_178_117_gat), .Y(G178_117_gat) );
BUFX20 U_g1166 (.A(GIN_179_118_gat), .Y(G179_118_gat) );
BUFX20 U_g1167 (.A(GIN_180_119_gat), .Y(G180_119_gat) );
BUFX20 U_g1168 (.A(GIN_181_120_gat), .Y(G181_120_gat) );
BUFX20 U_g1169 (.A(GIN_182_121_gat), .Y(G182_121_gat) );
BUFX20 U_g1170 (.A(GIN_183_122_gat), .Y(G183_122_gat) );
BUFX20 U_g1171 (.A(GIN_184_123_gat), .Y(G184_123_gat) );
BUFX20 U_g1172 (.A(GIN_185_124_gat), .Y(G185_124_gat) );
BUFX20 U_g1173 (.A(GIN_186_125_gat), .Y(G186_125_gat) );
BUFX20 U_g1174 (.A(GIN_189_126_gat), .Y(G189_126_gat) );
BUFX20 U_g1175 (.A(GIN_190_127_gat), .Y(G190_127_gat) );
BUFX20 U_g1176 (.A(GIN_191_128_gat), .Y(G191_128_gat) );
BUFX20 U_g1177 (.A(GIN_192_129_gat), .Y(G192_129_gat) );
BUFX20 U_g1178 (.A(GIN_193_130_gat), .Y(G193_130_gat) );
BUFX20 U_g1179 (.A(GIN_194_131_gat), .Y(G194_131_gat) );
BUFX20 U_g1180 (.A(GIN_195_132_gat), .Y(G195_132_gat) );
BUFX20 U_g1181 (.A(GIN_196_133_gat), .Y(G196_133_gat) );
BUFX20 U_g1182 (.A(GIN_197_134_gat), .Y(G197_134_gat) );
BUFX20 U_g1183 (.A(GIN_198_135_gat), .Y(G198_135_gat) );
BUFX20 U_g1184 (.A(GIN_199_136_gat), .Y(G199_136_gat) );
BUFX20 U_g1185 (.A(GIN_200_137_gat), .Y(G200_137_gat) );
BUFX20 U_g1186 (.A(GIN_201_138_gat), .Y(G201_138_gat) );
BUFX20 U_g1187 (.A(GIN_202_139_gat), .Y(G202_139_gat) );
BUFX20 U_g1188 (.A(GIN_203_140_gat), .Y(G203_140_gat) );
BUFX20 U_g1189 (.A(GIN_204_141_gat), .Y(G204_141_gat) );
BUFX20 U_g1190 (.A(GIN_205_142_gat), .Y(G205_142_gat) );
BUFX20 U_g1191 (.A(GIN_206_143_gat), .Y(G206_143_gat) );
BUFX20 U_g1192 (.A(GIN_207_144_gat), .Y(G207_144_gat) );
BUFX20 U_g1193 (.A(GIN_208_145_gat), .Y(G208_145_gat) );
BUFX20 U_g1194 (.A(GIN_209_146_gat), .Y(G209_146_gat) );
BUFX20 U_g1195 (.A(GIN_210_147_gat), .Y(G210_147_gat) );
BUFX20 U_g1196 (.A(GIN_211_148_gat), .Y(G211_148_gat) );
BUFX20 U_g1197 (.A(GIN_212_149_gat), .Y(G212_149_gat) );
BUFX20 U_g1198 (.A(GIN_213_150_gat), .Y(G213_150_gat) );
BUFX20 U_g1199 (.A(GIN_214_151_gat), .Y(G214_151_gat) );
BUFX20 U_g1200 (.A(GIN_215_152_gat), .Y(G215_152_gat) );
BUFX20 U_g1201 (.A(GIN_239_153_gat), .Y(G239_153_gat) );
BUFX20 U_g1202 (.A(GIN_240_154_gat), .Y(G240_154_gat) );
BUFX20 U_g1203 (.A(GIN_241_155_gat), .Y(G241_155_gat) );
BUFX20 U_g1204 (.A(GIN_242_156_gat), .Y(G242_156_gat) );
BUFX20 U_g1205 (.A(GIN_243_157_gat), .Y(G243_157_gat) );
BUFX20 U_g1206 (.A(GIN_244_158_gat), .Y(G244_158_gat) );
BUFX20 U_g1207 (.A(GIN_245_159_gat), .Y(G245_159_gat) );
BUFX20 U_g1208 (.A(GIN_246_160_gat), .Y(G246_160_gat) );
BUFX20 U_g1209 (.A(GIN_247_161_gat), .Y(G247_161_gat) );
BUFX20 U_g1210 (.A(GIN_248_162_gat), .Y(G248_162_gat) );
BUFX20 U_g1211 (.A(GIN_249_163_gat), .Y(G249_163_gat) );
BUFX20 U_g1212 (.A(GIN_250_164_gat), .Y(G250_164_gat) );
BUFX20 U_g1213 (.A(GIN_251_165_gat), .Y(G251_165_gat) );
BUFX20 U_g1214 (.A(GIN_252_166_gat), .Y(G252_166_gat) );
BUFX20 U_g1215 (.A(GIN_253_167_gat), .Y(G253_167_gat) );
BUFX20 U_g1216 (.A(GIN_254_168_gat), .Y(G254_168_gat) );
BUFX20 U_g1217 (.A(GIN_255_169_gat), .Y(G255_169_gat) );
BUFX20 U_g1218 (.A(GIN_256_170_gat), .Y(G256_170_gat) );
BUFX20 U_g1219 (.A(GIN_257_171_gat), .Y(G257_171_gat) );
BUFX20 U_g1220 (.A(GIN_262_172_gat), .Y(G262_172_gat) );
BUFX20 U_g1221 (.A(GIN_263_173_gat), .Y(G263_173_gat) );
BUFX20 U_g1222 (.A(GIN_264_174_gat), .Y(G264_174_gat) );
BUFX20 U_g1223 (.A(GIN_265_175_gat), .Y(G265_175_gat) );
BUFX20 U_g1224 (.A(GIN_266_176_gat), .Y(G266_176_gat) );
BUFX20 U_g1225 (.A(GIN_267_177_gat), .Y(G267_177_gat) );
BUFX20 U_g1226 (.A(GIN_268_178_gat), .Y(G268_178_gat) );
BUFX20 U_g1227 (.A(GIN_269_179_gat), .Y(G269_179_gat) );
BUFX20 U_g1228 (.A(GIN_270_180_gat), .Y(G270_180_gat) );
BUFX20 U_g1229 (.A(GIN_271_181_gat), .Y(G271_181_gat) );
BUFX20 U_g1230 (.A(GIN_272_182_gat), .Y(G272_182_gat) );
BUFX20 U_g1231 (.A(GIN_273_183_gat), .Y(G273_183_gat) );
BUFX20 U_g1232 (.A(GIN_274_184_gat), .Y(G274_184_gat) );
BUFX20 U_g1233 (.A(GIN_275_185_gat), .Y(G275_185_gat) );
BUFX20 U_g1234 (.A(GIN_276_186_gat), .Y(G276_186_gat) );
BUFX20 U_g1235 (.A(GIN_277_187_gat), .Y(G277_187_gat) );
BUFX20 U_g1236 (.A(GIN_278_188_gat), .Y(G278_188_gat) );
BUFX20 U_g1237 (.A(GIN_279_189_gat), .Y(G279_189_gat) );
BUFX20 U_g1238 (.A(G452_190_gat), .Y(G350_301_gat) );
BUFX20 U_g1239 (.A(G452_190_gat), .Y(G335_299_gat) );
BUFX20 U_g1240 (.A(G452_190_gat), .Y(G409_298_gat) );
BUFX20 U_g1241 (.A(G1083_199_gat), .Y(G369_289_gat) );
BUFX20 U_g1242 (.A(G1083_199_gat), .Y(G367_288_gat) );
BUFX20 U_g1243 (.A(G2066_212_gat), .Y(G411_264_gat) );
BUFX20 U_g1244 (.A(G2066_212_gat), .Y(G337_263_gat) );
BUFX20 U_g1245 (.A(G2066_212_gat), .Y(G384_262_gat) );
BUFX20 U_g1246 (.A(G897_755_gat), .Y(G284_847_gat) );
BUFX20 U_g1247 (.A(G897_755_gat), .Y(G321_848_gat) );
BUFX20 U_g1248 (.A(G898_756_gat), .Y(G297_849_gat) );
BUFX20 U_g1249 (.A(G898_756_gat), .Y(G280_850_gat) );
BUFX20 U_g1250 (.A(G896_846_gat), .Y(G282_922_gat) );
BUFX20 U_g1251 (.A(G896_846_gat), .Y(G323_923_gat) );
BUFX20 U_g1252 (.A(G895_1396_gat), .Y(G295_1400_gat) );
BUFX20 U_g1253 (.A(G895_1396_gat), .Y(G331_1401_gat) );
INVXL U_g1254 (.A(G567_194_gat), .Y(G567_194_ngat) );
INVXL U_g1255 (.A(G1955_320_gat), .Y(G1955_320_ngat) );
INVXL U_g1256 (.A(G154_964_gat), .Y(G154_964_ngat) );
INVXL U_g1257 (.A(G155_967_gat), .Y(G155_967_ngat) );
INVXL U_g1258 (.A(G2675_261_gat), .Y(G2675_261_ngat) );
INVXL U_g1259 (.A(G2682_233_gat), .Y(G2682_233_ngat) );
INVXL U_g1260 (.A(G2471_282_gat), .Y(G2471_282_ngat) );
INVXL U_g1261 (.A(G2478_234_gat), .Y(G2478_234_ngat) );
INVXL U_g1262 (.A(G2454_230_gat), .Y(G2454_230_ngat) );
INVXL U_g1263 (.A(G2457_236_gat), .Y(G2457_236_ngat) );
INVXL U_g1264 (.A(G2451_229_gat), .Y(G2451_229_ngat) );
INVXL U_g1265 (.A(G2458_235_gat), .Y(G2458_235_ngat) );
INVXL U_g1266 (.A(G2446_228_gat), .Y(G2446_228_ngat) );
INVXL U_g1267 (.A(G2449_238_gat), .Y(G2449_238_ngat) );
INVXL U_g1268 (.A(G2443_227_gat), .Y(G2443_227_ngat) );
INVXL U_g1269 (.A(G2450_237_gat), .Y(G2450_237_ngat) );
INVXL U_g1270 (.A(G2438_226_gat), .Y(G2438_226_ngat) );
INVXL U_g1271 (.A(G2441_240_gat), .Y(G2441_240_ngat) );
INVXL U_g1272 (.A(G2435_225_gat), .Y(G2435_225_ngat) );
INVXL U_g1273 (.A(G2442_239_gat), .Y(G2442_239_ngat) );
INVXL U_g1274 (.A(G2430_224_gat), .Y(G2430_224_ngat) );
INVXL U_g1275 (.A(G2433_242_gat), .Y(G2433_242_ngat) );
INVXL U_g1276 (.A(G2427_223_gat), .Y(G2427_223_ngat) );
INVXL U_g1277 (.A(G2434_241_gat), .Y(G2434_241_ngat) );
INVXL U_g1278 (.A(G2678_232_gat), .Y(G2678_232_ngat) );
INVXL U_g1279 (.A(G2681_351_gat), .Y(G2681_351_ngat) );
INVXL U_g1280 (.A(G2474_231_gat), .Y(G2474_231_ngat) );
INVXL U_g1281 (.A(G2477_369_gat), .Y(G2477_369_ngat) );
INVXL U_g1282 (.A(G2459_325_gat), .Y(G2459_325_ngat) );
INVXL U_g1283 (.A(G2460_326_gat), .Y(G2460_326_ngat) );
INVXL U_g1284 (.A(G1493_327_gat), .Y(G1493_327_ngat) );
INVXL U_g1285 (.A(G1494_328_gat), .Y(G1494_328_ngat) );
INVXL U_g1286 (.A(G1484_329_gat), .Y(G1484_329_ngat) );
INVXL U_g1287 (.A(G1485_330_gat), .Y(G1485_330_ngat) );
INVXL U_g1288 (.A(G1475_331_gat), .Y(G1475_331_ngat) );
INVXL U_g1289 (.A(G1476_332_gat), .Y(G1476_332_ngat) );
INVXL U_g1290 (.A(G2699_248_gat), .Y(G2699_248_ngat) );
INVXL U_g1291 (.A(G2706_340_gat), .Y(G2706_340_ngat) );
INVXL U_g1292 (.A(G2702_250_gat), .Y(G2702_250_ngat) );
INVXL U_g1293 (.A(G2705_339_gat), .Y(G2705_339_ngat) );
INVXL U_g1294 (.A(G2691_252_gat), .Y(G2691_252_ngat) );
INVXL U_g1295 (.A(G2698_344_gat), .Y(G2698_344_ngat) );
INVXL U_g1296 (.A(G2694_254_gat), .Y(G2694_254_ngat) );
INVXL U_g1297 (.A(G2697_342_gat), .Y(G2697_342_ngat) );
INVXL U_g1298 (.A(G2683_256_gat), .Y(G2683_256_ngat) );
INVXL U_g1299 (.A(G2690_348_gat), .Y(G2690_348_ngat) );
INVXL U_g1300 (.A(G2686_258_gat), .Y(G2686_258_ngat) );
INVXL U_g1301 (.A(G2689_346_gat), .Y(G2689_346_ngat) );
INVXL U_g1302 (.A(G2505_266_gat), .Y(G2505_266_ngat) );
INVXL U_g1303 (.A(G2512_355_gat), .Y(G2512_355_ngat) );
INVXL U_g1304 (.A(G2508_268_gat), .Y(G2508_268_ngat) );
INVXL U_g1305 (.A(G2511_353_gat), .Y(G2511_353_ngat) );
INVXL U_g1306 (.A(G2495_270_gat), .Y(G2495_270_ngat) );
INVXL U_g1307 (.A(G2502_359_gat), .Y(G2502_359_ngat) );
INVXL U_g1308 (.A(G2498_272_gat), .Y(G2498_272_ngat) );
INVXL U_g1309 (.A(G2501_357_gat), .Y(G2501_357_ngat) );
INVXL U_g1310 (.A(G2487_274_gat), .Y(G2487_274_ngat) );
INVXL U_g1311 (.A(G2494_363_gat), .Y(G2494_363_ngat) );
INVXL U_g1312 (.A(G2490_276_gat), .Y(G2490_276_ngat) );
INVXL U_g1313 (.A(G2493_361_gat), .Y(G2493_361_ngat) );
INVXL U_g1314 (.A(G2479_278_gat), .Y(G2479_278_ngat) );
INVXL U_g1315 (.A(G2486_367_gat), .Y(G2486_367_ngat) );
INVXL U_g1316 (.A(G2482_280_gat), .Y(G2482_280_ngat) );
INVXL U_g1317 (.A(G2485_365_gat), .Y(G2485_365_ngat) );
INVXL U_g1318 (.A(G2461_285_gat), .Y(G2461_285_ngat) );
INVXL U_g1319 (.A(G2468_373_gat), .Y(G2468_373_ngat) );
INVXL U_g1320 (.A(G2464_287_gat), .Y(G2464_287_ngat) );
INVXL U_g1321 (.A(G2467_371_gat), .Y(G2467_371_ngat) );
INVXL U_g1322 (.A(G1775_416_gat), .Y(G1775_416_ngat) );
INVXL U_g1323 (.A(G1776_323_gat), .Y(G1776_323_ngat) );
INVXL U_g1324 (.A(G1498_417_gat), .Y(G1498_417_ngat) );
INVXL U_g1325 (.A(G1499_324_gat), .Y(G1499_324_ngat) );
INVXL U_g1326 (.A(G2707_428_gat), .Y(G2707_428_ngat) );
INVXL U_g1327 (.A(G2708_427_gat), .Y(G2708_427_ngat) );
INVXL U_g1328 (.A(G1793_432_gat), .Y(G1793_432_ngat) );
INVXL U_g1329 (.A(G1794_430_gat), .Y(G1794_430_ngat) );
INVXL U_g1330 (.A(G1784_436_gat), .Y(G1784_436_ngat) );
INVXL U_g1331 (.A(G1785_434_gat), .Y(G1785_434_ngat) );
INVXL U_g1332 (.A(G2513_441_gat), .Y(G2513_441_ngat) );
INVXL U_g1333 (.A(G2514_439_gat), .Y(G2514_439_ngat) );
INVXL U_g1334 (.A(G2503_445_gat), .Y(G2503_445_ngat) );
INVXL U_g1335 (.A(G2504_443_gat), .Y(G2504_443_ngat) );
INVXL U_g1336 (.A(G1516_449_gat), .Y(G1516_449_ngat) );
INVXL U_g1337 (.A(G1517_447_gat), .Y(G1517_447_ngat) );
INVXL U_g1338 (.A(G1507_453_gat), .Y(G1507_453_ngat) );
INVXL U_g1339 (.A(G1508_451_gat), .Y(G1508_451_ngat) );
INVXL U_g1340 (.A(G2469_458_gat), .Y(G2469_458_ngat) );
INVXL U_g1341 (.A(G2470_456_gat), .Y(G2470_456_ngat) );
INVXL U_g1342 (.A(G2515_553_gat), .Y(G2515_553_ngat) );
INVXL U_g1343 (.A(G2522_539_gat), .Y(G2522_539_ngat) );
INVXL U_g1344 (.A(G2103_247_gat), .Y(G2103_247_ngat) );
INVXL U_g1345 (.A(G1473_545_gat), .Y(G1473_545_ngat) );
INVXL U_g1346 (.A(G2099_249_gat), .Y(G2099_249_ngat) );
INVXL U_g1347 (.A(G1470_562_gat), .Y(G1470_562_ngat) );
INVXL U_g1348 (.A(G2518_418_gat), .Y(G2518_418_ngat) );
INVXL U_g1349 (.A(G2521_595_gat), .Y(G2521_595_ngat) );
INVXL U_g1350 (.A(G2525_549_gat), .Y(G2525_549_ngat) );
INVXL U_g1351 (.A(G2532_590_gat), .Y(G2532_590_ngat) );
INVXL U_g1352 (.A(G2528_550_gat), .Y(G2528_550_ngat) );
INVXL U_g1353 (.A(G2531_589_gat), .Y(G2531_589_ngat) );
INVXL U_g1354 (.A(G560_295_gat), .Y(G560_295_ngat) );
INVXL U_g1355 (.A(G852_619_gat), .Y(G852_619_ngat) );
INVXL U_g1356 (.A(G2631_615_gat), .Y(G2631_615_ngat) );
INVXL U_g1357 (.A(G2638_602_gat), .Y(G2638_602_ngat) );
INVXL U_g1358 (.A(G2523_653_gat), .Y(G2523_653_ngat) );
INVXL U_g1359 (.A(G2524_576_gat), .Y(G2524_576_ngat) );
INVXL U_g1360 (.A(G1540_655_gat), .Y(G1540_655_ngat) );
INVXL U_g1361 (.A(G1541_577_gat), .Y(G1541_577_ngat) );
INVXL U_g1362 (.A(G1537_654_gat), .Y(G1537_654_ngat) );
INVXL U_g1363 (.A(G1538_580_gat), .Y(G1538_580_ngat) );
INVXL U_g1364 (.A(G2665_582_gat), .Y(G2665_582_ngat) );
INVXL U_g1365 (.A(G2672_682_gat), .Y(G2672_682_ngat) );
INVXL U_g1366 (.A(G2778_711_gat), .Y(G2778_711_ngat) );
INVXL U_g1367 (.A(G2781_429_gat), .Y(G2781_429_ngat) );
INVXL U_g1368 (.A(G2770_712_gat), .Y(G2770_712_ngat) );
INVXL U_g1369 (.A(G2773_431_gat), .Y(G2773_431_ngat) );
INVXL U_g1370 (.A(G2762_716_gat), .Y(G2762_716_ngat) );
INVXL U_g1371 (.A(G2765_433_gat), .Y(G2765_433_ngat) );
INVXL U_g1372 (.A(G2754_713_gat), .Y(G2754_713_ngat) );
INVXL U_g1373 (.A(G2757_435_gat), .Y(G2757_435_ngat) );
INVXL U_g1374 (.A(G2746_717_gat), .Y(G2746_717_ngat) );
INVXL U_g1375 (.A(G2749_437_gat), .Y(G2749_437_ngat) );
INVXL U_g1376 (.A(G2738_714_gat), .Y(G2738_714_ngat) );
INVXL U_g1377 (.A(G2741_438_gat), .Y(G2741_438_ngat) );
INVXL U_g1378 (.A(G2533_664_gat), .Y(G2533_664_ngat) );
INVXL U_g1379 (.A(G2534_663_gat), .Y(G2534_663_ngat) );
INVXL U_g1380 (.A(G2626_718_gat), .Y(G2626_718_ngat) );
INVXL U_g1381 (.A(G2629_440_gat), .Y(G2629_440_ngat) );
INVXL U_g1382 (.A(G2618_719_gat), .Y(G2618_719_ngat) );
INVXL U_g1383 (.A(G2621_442_gat), .Y(G2621_442_ngat) );
INVXL U_g1384 (.A(G2610_725_gat), .Y(G2610_725_ngat) );
INVXL U_g1385 (.A(G2613_444_gat), .Y(G2613_444_ngat) );
INVXL U_g1386 (.A(G2602_720_gat), .Y(G2602_720_ngat) );
INVXL U_g1387 (.A(G2605_446_gat), .Y(G2605_446_ngat) );
INVXL U_g1388 (.A(G2594_721_gat), .Y(G2594_721_ngat) );
INVXL U_g1389 (.A(G2597_448_gat), .Y(G2597_448_ngat) );
INVXL U_g1390 (.A(G2586_722_gat), .Y(G2586_722_ngat) );
INVXL U_g1391 (.A(G2589_450_gat), .Y(G2589_450_ngat) );
INVXL U_g1392 (.A(G2578_726_gat), .Y(G2578_726_ngat) );
INVXL U_g1393 (.A(G2581_452_gat), .Y(G2581_452_ngat) );
INVXL U_g1394 (.A(G2570_723_gat), .Y(G2570_723_ngat) );
INVXL U_g1395 (.A(G2573_454_gat), .Y(G2573_454_ngat) );
INVXL U_g1396 (.A(G2562_727_gat), .Y(G2562_727_ngat) );
INVXL U_g1397 (.A(G2565_455_gat), .Y(G2565_455_ngat) );
INVXL U_g1398 (.A(G2554_724_gat), .Y(G2554_724_ngat) );
INVXL U_g1399 (.A(G2557_457_gat), .Y(G2557_457_ngat) );
INVXL U_g1400 (.A(G2634_555_gat), .Y(G2634_555_ngat) );
INVXL U_g1401 (.A(G2637_683_gat), .Y(G2637_683_ngat) );
INVXL U_g1402 (.A(G2642_603_gat), .Y(G2642_603_ngat) );
INVXL U_g1403 (.A(G2645_676_gat), .Y(G2645_676_ngat) );
INVXL U_g1404 (.A(G2639_605_gat), .Y(G2639_605_ngat) );
INVXL U_g1405 (.A(G2646_675_gat), .Y(G2646_675_ngat) );
INVXL U_g1406 (.A(G2650_606_gat), .Y(G2650_606_ngat) );
INVXL U_g1407 (.A(G2653_678_gat), .Y(G2653_678_ngat) );
INVXL U_g1408 (.A(G2647_608_gat), .Y(G2647_608_ngat) );
INVXL U_g1409 (.A(G2654_677_gat), .Y(G2654_677_ngat) );
INVXL U_g1410 (.A(G2658_611_gat), .Y(G2658_611_ngat) );
INVXL U_g1411 (.A(G2661_680_gat), .Y(G2661_680_ngat) );
INVXL U_g1412 (.A(G2655_613_gat), .Y(G2655_613_ngat) );
INVXL U_g1413 (.A(G2662_679_gat), .Y(G2662_679_ngat) );
INVXL U_g1414 (.A(G2668_614_gat), .Y(G2668_614_ngat) );
INVXL U_g1415 (.A(G2671_658_gat), .Y(G2671_658_ngat) );
INVXL U_g1416 (.A(G2151_691_gat), .Y(G2151_691_ngat) );
INVXL U_g1417 (.A(G2158_708_gat), .Y(G2158_708_ngat) );
INVXL U_g1418 (.A(G1820_739_gat), .Y(G1820_739_ngat) );
INVXL U_g1419 (.A(G1821_649_gat), .Y(G1821_649_ngat) );
INVXL U_g1420 (.A(G1823_728_gat), .Y(G1823_728_ngat) );
INVXL U_g1421 (.A(G1824_650_gat), .Y(G1824_650_ngat) );
INVXL U_g1422 (.A(G1543_750_gat), .Y(G1543_750_ngat) );
INVXL U_g1423 (.A(G1544_651_gat), .Y(G1544_651_ngat) );
INVXL U_g1424 (.A(G1546_729_gat), .Y(G1546_729_ngat) );
INVXL U_g1425 (.A(G1547_652_gat), .Y(G1547_652_ngat) );
INVXL U_g1426 (.A(G1542_731_gat), .Y(G1542_731_ngat) );
INVXL U_g1427 (.A(G1539_732_gat), .Y(G1539_732_ngat) );
INVXL U_g1428 (.A(G2673_769_gat), .Y(G2673_769_ngat) );
INVXL U_g1429 (.A(G2674_734_gat), .Y(G2674_734_ngat) );
INVXL U_g1430 (.A(G2775_341_gat), .Y(G2775_341_ngat) );
INVXL U_g1431 (.A(G2782_804_gat), .Y(G2782_804_ngat) );
INVXL U_g1432 (.A(G2767_343_gat), .Y(G2767_343_ngat) );
INVXL U_g1433 (.A(G2774_805_gat), .Y(G2774_805_ngat) );
INVXL U_g1434 (.A(G2759_345_gat), .Y(G2759_345_ngat) );
INVXL U_g1435 (.A(G2766_808_gat), .Y(G2766_808_ngat) );
INVXL U_g1436 (.A(G2751_347_gat), .Y(G2751_347_ngat) );
INVXL U_g1437 (.A(G2758_806_gat), .Y(G2758_806_ngat) );
INVXL U_g1438 (.A(G2743_350_gat), .Y(G2743_350_ngat) );
INVXL U_g1439 (.A(G2750_809_gat), .Y(G2750_809_ngat) );
INVXL U_g1440 (.A(G2735_352_gat), .Y(G2735_352_ngat) );
INVXL U_g1441 (.A(G2742_807_gat), .Y(G2742_807_ngat) );
INVXL U_g1442 (.A(G2623_354_gat), .Y(G2623_354_ngat) );
INVXL U_g1443 (.A(G2630_810_gat), .Y(G2630_810_ngat) );
INVXL U_g1444 (.A(G2615_356_gat), .Y(G2615_356_ngat) );
INVXL U_g1445 (.A(G2622_811_gat), .Y(G2622_811_ngat) );
INVXL U_g1446 (.A(G2607_358_gat), .Y(G2607_358_ngat) );
INVXL U_g1447 (.A(G2614_817_gat), .Y(G2614_817_ngat) );
INVXL U_g1448 (.A(G2599_360_gat), .Y(G2599_360_ngat) );
INVXL U_g1449 (.A(G2606_812_gat), .Y(G2606_812_ngat) );
INVXL U_g1450 (.A(G2591_362_gat), .Y(G2591_362_ngat) );
INVXL U_g1451 (.A(G2598_813_gat), .Y(G2598_813_ngat) );
INVXL U_g1452 (.A(G2583_364_gat), .Y(G2583_364_ngat) );
INVXL U_g1453 (.A(G2590_814_gat), .Y(G2590_814_ngat) );
INVXL U_g1454 (.A(G2575_366_gat), .Y(G2575_366_ngat) );
INVXL U_g1455 (.A(G2582_818_gat), .Y(G2582_818_ngat) );
INVXL U_g1456 (.A(G2567_368_gat), .Y(G2567_368_ngat) );
INVXL U_g1457 (.A(G2574_815_gat), .Y(G2574_815_ngat) );
INVXL U_g1458 (.A(G2559_370_gat), .Y(G2559_370_ngat) );
INVXL U_g1459 (.A(G2566_819_gat), .Y(G2566_819_ngat) );
INVXL U_g1460 (.A(G2551_372_gat), .Y(G2551_372_ngat) );
INVXL U_g1461 (.A(G2558_816_gat), .Y(G2558_816_ngat) );
INVXL U_g1462 (.A(G1752_762_gat), .Y(G1752_762_ngat) );
INVXL U_g1463 (.A(G1753_674_gat), .Y(G1753_674_ngat) );
INVXL U_g1464 (.A(G1761_763_gat), .Y(G1761_763_ngat) );
INVXL U_g1465 (.A(G1762_764_gat), .Y(G1762_764_ngat) );
INVXL U_g1466 (.A(G1770_765_gat), .Y(G1770_765_ngat) );
INVXL U_g1467 (.A(G1771_766_gat), .Y(G1771_766_ngat) );
INVXL U_g1468 (.A(G2663_767_gat), .Y(G2663_767_ngat) );
INVXL U_g1469 (.A(G2664_768_gat), .Y(G2664_768_ngat) );
INVXL U_g1470 (.A(G2110_685_gat), .Y(G2110_685_ngat) );
INVXL U_g1471 (.A(G2113_795_gat), .Y(G2113_795_ngat) );
INVXL U_g1472 (.A(G2164_686_gat), .Y(G2164_686_ngat) );
INVXL U_g1473 (.A(G2167_796_gat), .Y(G2167_796_ngat) );
INVXL U_g1474 (.A(G2115_780_gat), .Y(G2115_780_ngat) );
INVXL U_g1475 (.A(G2122_774_gat), .Y(G2122_774_ngat) );
INVXL U_g1476 (.A(G2169_782_gat), .Y(G2169_782_ngat) );
INVXL U_g1477 (.A(G2176_776_gat), .Y(G2176_776_ngat) );
INVXL U_g1478 (.A(G2126_785_gat), .Y(G2126_785_ngat) );
INVXL U_g1479 (.A(G2129_786_gat), .Y(G2129_786_ngat) );
INVXL U_g1480 (.A(G2107_706_gat), .Y(G2107_706_ngat) );
INVXL U_g1481 (.A(G2114_771_gat), .Y(G2114_771_ngat) );
INVXL U_g1482 (.A(G2161_707_gat), .Y(G2161_707_ngat) );
INVXL U_g1483 (.A(G2168_772_gat), .Y(G2168_772_ngat) );
INVXL U_g1484 (.A(G2154_631_gat), .Y(G2154_631_ngat) );
INVXL U_g1485 (.A(G2157_777_gat), .Y(G2157_777_ngat) );
INVXL U_g1486 (.A(G1825_821_gat), .Y(G1825_821_ngat) );
INVXL U_g1487 (.A(G1822_820_gat), .Y(G1822_820_ngat) );
INVXL U_g1488 (.A(G1548_823_gat), .Y(G1548_823_ngat) );
INVXL U_g1489 (.A(G1545_822_gat), .Y(G1545_822_ngat) );
INVXL U_g1490 (.A(G2535_825_gat), .Y(G2535_825_ngat) );
INVXL U_g1491 (.A(G2542_824_gat), .Y(G2542_824_ngat) );
INVXL U_g1492 (.A(G2059_736_gat), .Y(G2059_736_ngat) );
INVXL U_g1493 (.A(G2060_829_gat), .Y(G2060_829_ngat) );
INVXL U_g1494 (.A(G2055_737_gat), .Y(G2055_737_ngat) );
INVXL U_g1495 (.A(G2056_830_gat), .Y(G2056_830_ngat) );
INVXL U_g1496 (.A(G2051_738_gat), .Y(G2051_738_ngat) );
INVXL U_g1497 (.A(G2052_831_gat), .Y(G2052_831_ngat) );
INVXL U_g1498 (.A(G2047_740_gat), .Y(G2047_740_ngat) );
INVXL U_g1499 (.A(G2048_832_gat), .Y(G2048_832_ngat) );
INVXL U_g1500 (.A(G2043_741_gat), .Y(G2043_741_ngat) );
INVXL U_g1501 (.A(G2044_833_gat), .Y(G2044_833_ngat) );
INVXL U_g1502 (.A(G2039_742_gat), .Y(G2039_742_ngat) );
INVXL U_g1503 (.A(G2040_834_gat), .Y(G2040_834_ngat) );
INVXL U_g1504 (.A(G1597_744_gat), .Y(G1597_744_ngat) );
INVXL U_g1505 (.A(G1598_836_gat), .Y(G1598_836_ngat) );
INVXL U_g1506 (.A(G1593_745_gat), .Y(G1593_745_ngat) );
INVXL U_g1507 (.A(G1594_837_gat), .Y(G1594_837_ngat) );
INVXL U_g1508 (.A(G1589_746_gat), .Y(G1589_746_ngat) );
INVXL U_g1509 (.A(G1590_838_gat), .Y(G1590_838_ngat) );
INVXL U_g1510 (.A(G1585_747_gat), .Y(G1585_747_ngat) );
INVXL U_g1511 (.A(G1586_839_gat), .Y(G1586_839_ngat) );
INVXL U_g1512 (.A(G1581_748_gat), .Y(G1581_748_ngat) );
INVXL U_g1513 (.A(G1582_840_gat), .Y(G1582_840_ngat) );
INVXL U_g1514 (.A(G1577_749_gat), .Y(G1577_749_ngat) );
INVXL U_g1515 (.A(G1578_841_gat), .Y(G1578_841_ngat) );
INVXL U_g1516 (.A(G1573_751_gat), .Y(G1573_751_ngat) );
INVXL U_g1517 (.A(G1574_842_gat), .Y(G1574_842_ngat) );
INVXL U_g1518 (.A(G1569_752_gat), .Y(G1569_752_ngat) );
INVXL U_g1519 (.A(G1570_843_gat), .Y(G1570_843_ngat) );
INVXL U_g1520 (.A(G1565_753_gat), .Y(G1565_753_ngat) );
INVXL U_g1521 (.A(G1566_844_gat), .Y(G1566_844_ngat) );
INVXL U_g1522 (.A(G1561_754_gat), .Y(G1561_754_ngat) );
INVXL U_g1523 (.A(G1562_845_gat), .Y(G1562_845_ngat) );
INVXL U_g1524 (.A(G569_864_gat), .Y(G569_864_ngat) );
INVXL U_g1525 (.A(G570_890_gat), .Y(G570_890_ngat) );
INVXL U_g1526 (.A(G599_865_gat), .Y(G599_865_ngat) );
INVXL U_g1527 (.A(G600_891_gat), .Y(G600_891_ngat) );
INVXL U_g1528 (.A(G2118_688_gat), .Y(G2118_688_ngat) );
INVXL U_g1529 (.A(G2121_869_gat), .Y(G2121_869_ngat) );
INVXL U_g1530 (.A(G2172_690_gat), .Y(G2172_690_ngat) );
INVXL U_g1531 (.A(G2175_871_gat), .Y(G2175_871_ngat) );
INVXL U_g1532 (.A(G2159_892_gat), .Y(G2159_892_ngat) );
INVXL U_g1533 (.A(G2160_778_gat), .Y(G2160_778_ngat) );
INVXL U_g1534 (.A(G2123_697_gat), .Y(G2123_697_ngat) );
INVXL U_g1535 (.A(G2130_875_gat), .Y(G2130_875_ngat) );
INVXL U_g1536 (.A(G2134_787_gat), .Y(G2134_787_ngat) );
INVXL U_g1537 (.A(G2137_882_gat), .Y(G2137_882_ngat) );
INVXL U_g1538 (.A(G2180_788_gat), .Y(G2180_788_ngat) );
INVXL U_g1539 (.A(G2183_883_gat), .Y(G2183_883_ngat) );
INVXL U_g1540 (.A(G2131_789_gat), .Y(G2131_789_ngat) );
INVXL U_g1541 (.A(G2138_880_gat), .Y(G2138_880_ngat) );
INVXL U_g1542 (.A(G2177_790_gat), .Y(G2177_790_ngat) );
INVXL U_g1543 (.A(G2184_881_gat), .Y(G2184_881_ngat) );
INVXL U_g1544 (.A(G2144_791_gat), .Y(G2144_791_ngat) );
INVXL U_g1545 (.A(G2147_888_gat), .Y(G2147_888_ngat) );
INVXL U_g1546 (.A(G2190_792_gat), .Y(G2190_792_ngat) );
INVXL U_g1547 (.A(G2193_889_gat), .Y(G2193_889_ngat) );
INVXL U_g1548 (.A(G2141_793_gat), .Y(G2141_793_ngat) );
INVXL U_g1549 (.A(G2148_884_gat), .Y(G2148_884_ngat) );
INVXL U_g1550 (.A(G2187_794_gat), .Y(G2187_794_ngat) );
INVXL U_g1551 (.A(G2194_885_gat), .Y(G2194_885_ngat) );
INVXL U_g1552 (.A(G2538_730_gat), .Y(G2538_730_ngat) );
INVXL U_g1553 (.A(G2541_902_gat), .Y(G2541_902_ngat) );
INVXL U_g1554 (.A(G2709_827_gat), .Y(G2709_827_ngat) );
INVXL U_g1555 (.A(G2716_928_gat), .Y(G2716_928_ngat) );
INVXL U_g1556 (.A(G2727_899_gat), .Y(G2727_899_ngat) );
INVXL U_g1557 (.A(G2734_584_gat), .Y(G2734_584_ngat) );
INVXL U_g1558 (.A(G2543_900_gat), .Y(G2543_900_ngat) );
INVXL U_g1559 (.A(G2550_835_gat), .Y(G2550_835_ngat) );
INVXL U_g1560 (.A(G2210_933_gat), .Y(G2210_933_ngat) );
INVXL U_g1561 (.A(G2213_852_gat), .Y(G2213_852_ngat) );
INVXL U_g1562 (.A(G2712_861_gat), .Y(G2712_861_ngat) );
INVXL U_g1563 (.A(G2715_904_gat), .Y(G2715_904_ngat) );
INVXL U_g1564 (.A(G578_931_gat), .Y(G578_931_ngat) );
INVXL U_g1565 (.A(G579_866_gat), .Y(G579_866_ngat) );
INVXL U_g1566 (.A(G608_932_gat), .Y(G608_932_ngat) );
INVXL U_g1567 (.A(G609_867_gat), .Y(G609_867_ngat) );
INVXL U_g1568 (.A(G587_874_gat), .Y(G587_874_ngat) );
INVXL U_g1569 (.A(G588_936_gat), .Y(G588_936_ngat) );
INVXL U_g1570 (.A(G2139_939_gat), .Y(G2139_939_ngat) );
INVXL U_g1571 (.A(G2140_943_gat), .Y(G2140_943_ngat) );
INVXL U_g1572 (.A(G2185_940_gat), .Y(G2185_940_ngat) );
INVXL U_g1573 (.A(G2186_944_gat), .Y(G2186_944_ngat) );
INVXL U_g1574 (.A(G2149_947_gat), .Y(G2149_947_ngat) );
INVXL U_g1575 (.A(G2150_949_gat), .Y(G2150_949_ngat) );
INVXL U_g1576 (.A(G2195_948_gat), .Y(G2195_948_ngat) );
INVXL U_g1577 (.A(G2196_950_gat), .Y(G2196_950_ngat) );
INVXL U_g1578 (.A(G1549_963_gat), .Y(G1549_963_ngat) );
INVXL U_g1579 (.A(G1550_901_gat), .Y(G1550_901_ngat) );
INVXL U_g1580 (.A(G2717_1018_gat), .Y(G2717_1018_ngat) );
INVXL U_g1581 (.A(G2718_965_gat), .Y(G2718_965_ngat) );
INVXL U_g1582 (.A(G2730_546_gat), .Y(G2730_546_ngat) );
INVXL U_g1583 (.A(G2733_961_gat), .Y(G2733_961_ngat) );
INVXL U_g1584 (.A(G2546_743_gat), .Y(G2546_743_ngat) );
INVXL U_g1585 (.A(G2549_962_gat), .Y(G2549_962_ngat) );
INVXL U_g1586 (.A(G2207_759_gat), .Y(G2207_759_ngat) );
INVXL U_g1587 (.A(G2214_1025_gat), .Y(G2214_1025_ngat) );
INVXL U_g1588 (.A(G1828_1048_gat), .Y(G1828_1048_ngat) );
INVXL U_g1589 (.A(G1829_966_gat), .Y(G1829_966_ngat) );
INVXL U_g1590 (.A(G1551_1062_gat), .Y(G1551_1062_ngat) );
INVXL U_g1591 (.A(G1552_978_gat), .Y(G1552_978_ngat) );
INVXL U_g1592 (.A(G2215_1009_gat), .Y(G2215_1009_ngat) );
INVXL U_g1593 (.A(G2216_1065_gat), .Y(G2216_1065_ngat) );
INVXL U_g1594 (.A(G1814_1069_gat), .Y(G1814_1069_ngat) );
INVXL U_g1595 (.A(G1815_1010_gat), .Y(G1815_1010_ngat) );
INVXL U_g1596 (.A(G1817_1066_gat), .Y(G1817_1066_ngat) );
INVXL U_g1597 (.A(G1818_1011_gat), .Y(G1818_1011_ngat) );
INVXL U_g1598 (.A(G2200_1031_gat), .Y(G2200_1031_ngat) );
INVXL U_g1599 (.A(G2203_1081_gat), .Y(G2203_1081_ngat) );
INVXL U_g1600 (.A(G2220_1032_gat), .Y(G2220_1032_ngat) );
INVXL U_g1601 (.A(G2223_1082_gat), .Y(G2223_1082_ngat) );
INVXL U_g1602 (.A(G2197_1033_gat), .Y(G2197_1033_ngat) );
INVXL U_g1603 (.A(G2204_1079_gat), .Y(G2204_1079_ngat) );
INVXL U_g1604 (.A(G2217_1034_gat), .Y(G2217_1034_ngat) );
INVXL U_g1605 (.A(G2224_1080_gat), .Y(G2224_1080_ngat) );
INVXL U_g1606 (.A(G1819_1128_gat), .Y(G1819_1128_ngat) );
INVXL U_g1607 (.A(G1816_1127_gat), .Y(G1816_1127_ngat) );
INVXL U_g1608 (.A(G2238_1124_gat), .Y(G2238_1124_ngat) );
INVXL U_g1609 (.A(G2241_770_gat), .Y(G2241_770_ngat) );
INVXL U_g1610 (.A(G2205_1147_gat), .Y(G2205_1147_ngat) );
INVXL U_g1611 (.A(G2206_1149_gat), .Y(G2206_1149_ngat) );
INVXL U_g1612 (.A(G2225_1148_gat), .Y(G2225_1148_ngat) );
INVXL U_g1613 (.A(G2226_1150_gat), .Y(G2226_1150_ngat) );
INVXL U_g1614 (.A(G2719_1190_gat), .Y(G2719_1190_ngat) );
INVXL U_g1615 (.A(G2726_1107_gat), .Y(G2726_1107_ngat) );
INVXL U_g1616 (.A(G635_1189_gat), .Y(G635_1189_ngat) );
INVXL U_g1617 (.A(G636_1125_gat), .Y(G636_1125_ngat) );
INVXL U_g1618 (.A(G638_1188_gat), .Y(G638_1188_ngat) );
INVXL U_g1619 (.A(G639_1126_gat), .Y(G639_1126_ngat) );
INVXL U_g1620 (.A(G2278_1130_gat), .Y(G2278_1130_ngat) );
INVXL U_g1621 (.A(G2281_1212_gat), .Y(G2281_1212_ngat) );
INVXL U_g1622 (.A(G2366_1132_gat), .Y(G2366_1132_ngat) );
INVXL U_g1623 (.A(G2369_1216_gat), .Y(G2369_1216_ngat) );
INVXL U_g1624 (.A(G2270_1134_gat), .Y(G2270_1134_ngat) );
INVXL U_g1625 (.A(G2273_1215_gat), .Y(G2273_1215_ngat) );
INVXL U_g1626 (.A(G2358_1136_gat), .Y(G2358_1136_ngat) );
INVXL U_g1627 (.A(G2361_1219_gat), .Y(G2361_1219_ngat) );
INVXL U_g1628 (.A(G2286_1138_gat), .Y(G2286_1138_ngat) );
INVXL U_g1629 (.A(G2289_1213_gat), .Y(G2289_1213_ngat) );
INVXL U_g1630 (.A(G2374_1140_gat), .Y(G2374_1140_ngat) );
INVXL U_g1631 (.A(G2377_1217_gat), .Y(G2377_1217_ngat) );
INVXL U_g1632 (.A(G2235_684_gat), .Y(G2235_684_ngat) );
INVXL U_g1633 (.A(G2242_1187_gat), .Y(G2242_1187_ngat) );
INVXL U_g1634 (.A(G629_1199_gat), .Y(G629_1199_ngat) );
INVXL U_g1635 (.A(G630_1141_gat), .Y(G630_1141_ngat) );
INVXL U_g1636 (.A(G632_1198_gat), .Y(G632_1198_ngat) );
INVXL U_g1637 (.A(G633_1142_gat), .Y(G633_1142_ngat) );
INVXL U_g1638 (.A(G2347_1185_gat), .Y(G2347_1185_ngat) );
INVXL U_g1639 (.A(G2354_773_gat), .Y(G2354_773_ngat) );
INVXL U_g1640 (.A(G2259_1186_gat), .Y(G2259_1186_ngat) );
INVXL U_g1641 (.A(G2266_775_gat), .Y(G2266_775_ngat) );
INVXL U_g1642 (.A(G2339_1184_gat), .Y(G2339_1184_ngat) );
INVXL U_g1643 (.A(G2346_868_gat), .Y(G2346_868_ngat) );
INVXL U_g1644 (.A(G2251_1183_gat), .Y(G2251_1183_ngat) );
INVXL U_g1645 (.A(G2258_870_gat), .Y(G2258_870_ngat) );
INVXL U_g1646 (.A(G2419_1182_gat), .Y(G2419_1182_ngat) );
INVXL U_g1647 (.A(G2426_872_gat), .Y(G2426_872_ngat) );
INVXL U_g1648 (.A(G2331_1181_gat), .Y(G2331_1181_ngat) );
INVXL U_g1649 (.A(G2338_873_gat), .Y(G2338_873_ngat) );
INVXL U_g1650 (.A(G2294_1152_gat), .Y(G2294_1152_ngat) );
INVXL U_g1651 (.A(G2297_1214_gat), .Y(G2297_1214_ngat) );
INVXL U_g1652 (.A(G2382_1154_gat), .Y(G2382_1154_ngat) );
INVXL U_g1653 (.A(G2385_1218_gat), .Y(G2385_1218_ngat) );
INVXL U_g1654 (.A(G2275_1155_gat), .Y(G2275_1155_ngat) );
INVXL U_g1655 (.A(G2282_1191_gat), .Y(G2282_1191_ngat) );
INVXL U_g1656 (.A(G2283_1156_gat), .Y(G2283_1156_ngat) );
INVXL U_g1657 (.A(G2290_1195_gat), .Y(G2290_1195_ngat) );
INVXL U_g1658 (.A(G2291_1157_gat), .Y(G2291_1157_ngat) );
INVXL U_g1659 (.A(G2298_1208_gat), .Y(G2298_1208_ngat) );
INVXL U_g1660 (.A(G2267_1158_gat), .Y(G2267_1158_ngat) );
INVXL U_g1661 (.A(G2274_1193_gat), .Y(G2274_1193_ngat) );
INVXL U_g1662 (.A(G2363_1159_gat), .Y(G2363_1159_ngat) );
INVXL U_g1663 (.A(G2370_1192_gat), .Y(G2370_1192_ngat) );
INVXL U_g1664 (.A(G2371_1160_gat), .Y(G2371_1160_ngat) );
INVXL U_g1665 (.A(G2378_1196_gat), .Y(G2378_1196_ngat) );
INVXL U_g1666 (.A(G2379_1161_gat), .Y(G2379_1161_ngat) );
INVXL U_g1667 (.A(G2386_1209_gat), .Y(G2386_1209_ngat) );
INVXL U_g1668 (.A(G2355_1162_gat), .Y(G2355_1162_ngat) );
INVXL U_g1669 (.A(G2362_1194_gat), .Y(G2362_1194_ngat) );
INVXL U_g1670 (.A(G2299_1164_gat), .Y(G2299_1164_ngat) );
INVXL U_g1671 (.A(G2306_1233_gat), .Y(G2306_1233_ngat) );
INVXL U_g1672 (.A(G2307_1166_gat), .Y(G2307_1166_ngat) );
INVXL U_g1673 (.A(G2314_1232_gat), .Y(G2314_1232_ngat) );
INVXL U_g1674 (.A(G2387_1168_gat), .Y(G2387_1168_ngat) );
INVXL U_g1675 (.A(G2394_1237_gat), .Y(G2394_1237_ngat) );
INVXL U_g1676 (.A(G2395_1170_gat), .Y(G2395_1170_ngat) );
INVXL U_g1677 (.A(G2402_1236_gat), .Y(G2402_1236_ngat) );
INVXL U_g1678 (.A(G2310_1173_gat), .Y(G2310_1173_ngat) );
INVXL U_g1679 (.A(G2313_1223_gat), .Y(G2313_1223_ngat) );
INVXL U_g1680 (.A(G2302_1174_gat), .Y(G2302_1174_ngat) );
INVXL U_g1681 (.A(G2305_1222_gat), .Y(G2305_1222_ngat) );
INVXL U_g1682 (.A(G2398_1177_gat), .Y(G2398_1177_ngat) );
INVXL U_g1683 (.A(G2401_1227_gat), .Y(G2401_1227_ngat) );
INVXL U_g1684 (.A(G2390_1178_gat), .Y(G2390_1178_ngat) );
INVXL U_g1685 (.A(G2393_1226_gat), .Y(G2393_1226_ngat) );
INVXL U_g1686 (.A(G2722_1047_gat), .Y(G2722_1047_ngat) );
INVXL U_g1687 (.A(G2725_1247_gat), .Y(G2725_1247_ngat) );
INVXL U_g1688 (.A(G640_1246_gat), .Y(G640_1246_ngat) );
INVXL U_g1689 (.A(G637_1245_gat), .Y(G637_1245_ngat) );
INVXL U_g1690 (.A(G908_1248_gat), .Y(G908_1248_ngat) );
INVXL U_g1691 (.A(G909_1267_gat), .Y(G909_1267_ngat) );
INVXL U_g1692 (.A(G1126_1249_gat), .Y(G1126_1249_ngat) );
INVXL U_g1693 (.A(G1127_1271_gat), .Y(G1127_1271_ngat) );
INVXL U_g1694 (.A(G899_1250_gat), .Y(G899_1250_ngat) );
INVXL U_g1695 (.A(G900_1270_gat), .Y(G900_1270_ngat) );
INVXL U_g1696 (.A(G1117_1251_gat), .Y(G1117_1251_ngat) );
INVXL U_g1697 (.A(G1118_1274_gat), .Y(G1118_1274_ngat) );
INVXL U_g1698 (.A(G916_1252_gat), .Y(G916_1252_ngat) );
INVXL U_g1699 (.A(G917_1268_gat), .Y(G917_1268_ngat) );
INVXL U_g1700 (.A(G1134_1253_gat), .Y(G1134_1253_ngat) );
INVXL U_g1701 (.A(G1135_1272_gat), .Y(G1135_1272_ngat) );
INVXL U_g1702 (.A(G645_1197_gat), .Y(G645_1197_ngat) );
INVXL U_g1703 (.A(G646_1254_gat), .Y(G646_1254_ngat) );
INVXL U_g1704 (.A(G634_1256_gat), .Y(G634_1256_ngat) );
INVXL U_g1705 (.A(G631_1255_gat), .Y(G631_1255_ngat) );
INVXL U_g1706 (.A(G2350_687_gat), .Y(G2350_687_ngat) );
INVXL U_g1707 (.A(G2353_1243_gat), .Y(G2353_1243_ngat) );
INVXL U_g1708 (.A(G2262_689_gat), .Y(G2262_689_ngat) );
INVXL U_g1709 (.A(G2265_1244_gat), .Y(G2265_1244_ngat) );
INVXL U_g1710 (.A(G2342_779_gat), .Y(G2342_779_ngat) );
INVXL U_g1711 (.A(G2345_1242_gat), .Y(G2345_1242_ngat) );
INVXL U_g1712 (.A(G2254_781_gat), .Y(G2254_781_ngat) );
INVXL U_g1713 (.A(G2257_1241_gat), .Y(G2257_1241_ngat) );
INVXL U_g1714 (.A(G2422_783_gat), .Y(G2422_783_ngat) );
INVXL U_g1715 (.A(G2425_1240_gat), .Y(G2425_1240_ngat) );
INVXL U_g1716 (.A(G2334_784_gat), .Y(G2334_784_ngat) );
INVXL U_g1717 (.A(G2337_1239_gat), .Y(G2337_1239_ngat) );
INVXL U_g1718 (.A(G925_1265_gat), .Y(G925_1265_ngat) );
INVXL U_g1719 (.A(G926_1269_gat), .Y(G926_1269_ngat) );
INVXL U_g1720 (.A(G1143_1266_gat), .Y(G1143_1266_ngat) );
INVXL U_g1721 (.A(G1144_1273_gat), .Y(G1144_1273_ngat) );
INVXL U_g1722 (.A(G928_1292_gat), .Y(G928_1292_ngat) );
INVXL U_g1723 (.A(G929_1279_gat), .Y(G929_1279_ngat) );
INVXL U_g1724 (.A(G938_1291_gat), .Y(G938_1291_ngat) );
INVXL U_g1725 (.A(G939_1280_gat), .Y(G939_1280_ngat) );
INVXL U_g1726 (.A(G2315_1281_gat), .Y(G2315_1281_ngat) );
INVXL U_g1727 (.A(G2322_1290_gat), .Y(G2322_1290_ngat) );
INVXL U_g1728 (.A(G2323_1282_gat), .Y(G2323_1282_ngat) );
INVXL U_g1729 (.A(G2330_1287_gat), .Y(G2330_1287_ngat) );
INVXL U_g1730 (.A(G1146_1298_gat), .Y(G1146_1298_ngat) );
INVXL U_g1731 (.A(G1147_1283_gat), .Y(G1147_1283_ngat) );
INVXL U_g1732 (.A(G1156_1297_gat), .Y(G1156_1297_ngat) );
INVXL U_g1733 (.A(G1157_1284_gat), .Y(G1157_1284_ngat) );
INVXL U_g1734 (.A(G2403_1285_gat), .Y(G2403_1285_ngat) );
INVXL U_g1735 (.A(G2410_1296_gat), .Y(G2410_1296_ngat) );
INVXL U_g1736 (.A(G2411_1286_gat), .Y(G2411_1286_ngat) );
INVXL U_g1737 (.A(G2418_1293_gat), .Y(G2418_1293_ngat) );
INVXL U_g1738 (.A(G1826_1299_gat), .Y(G1826_1299_ngat) );
INVXL U_g1739 (.A(G1827_1238_gat), .Y(G1827_1238_ngat) );
INVXL U_g1740 (.A(G1114_1309_gat), .Y(G1114_1309_ngat) );
INVXL U_g1741 (.A(G1115_1257_gat), .Y(G1115_1257_ngat) );
INVXL U_g1742 (.A(G683_1310_gat), .Y(G683_1310_ngat) );
INVXL U_g1743 (.A(G684_1258_gat), .Y(G684_1258_ngat) );
INVXL U_g1744 (.A(G1098_1311_gat), .Y(G1098_1311_ngat) );
INVXL U_g1745 (.A(G1099_1259_gat), .Y(G1099_1259_ngat) );
INVXL U_g1746 (.A(G664_1312_gat), .Y(G664_1312_ngat) );
INVXL U_g1747 (.A(G665_1260_gat), .Y(G665_1260_ngat) );
INVXL U_g1748 (.A(G1180_1313_gat), .Y(G1180_1313_ngat) );
INVXL U_g1749 (.A(G1181_1261_gat), .Y(G1181_1261_ngat) );
INVXL U_g1750 (.A(G962_1314_gat), .Y(G962_1314_ngat) );
INVXL U_g1751 (.A(G963_1262_gat), .Y(G963_1262_ngat) );
INVXL U_g1752 (.A(G2227_1308_gat), .Y(G2227_1308_ngat) );
INVXL U_g1753 (.A(G2234_1263_gat), .Y(G2234_1263_ngat) );
INVXL U_g1754 (.A(G2243_1300_gat), .Y(G2243_1300_ngat) );
INVXL U_g1755 (.A(G2250_1264_gat), .Y(G2250_1264_ngat) );
INVXL U_g1756 (.A(G2326_1230_gat), .Y(G2326_1230_ngat) );
INVXL U_g1757 (.A(G2329_1322_gat), .Y(G2329_1322_ngat) );
INVXL U_g1758 (.A(G2318_1231_gat), .Y(G2318_1231_ngat) );
INVXL U_g1759 (.A(G2321_1320_gat), .Y(G2321_1320_ngat) );
INVXL U_g1760 (.A(G2414_1234_gat), .Y(G2414_1234_ngat) );
INVXL U_g1761 (.A(G2417_1328_gat), .Y(G2417_1328_ngat) );
INVXL U_g1762 (.A(G2406_1235_gat), .Y(G2406_1235_ngat) );
INVXL U_g1763 (.A(G2409_1326_gat), .Y(G2409_1326_ngat) );
INVXL U_g1764 (.A(G2230_1206_gat), .Y(G2230_1206_ngat) );
INVXL U_g1765 (.A(G2233_1338_gat), .Y(G2233_1338_ngat) );
INVXL U_g1766 (.A(G2246_1207_gat), .Y(G2246_1207_ngat) );
INVXL U_g1767 (.A(G2249_1331_gat), .Y(G2249_1331_ngat) );
INVXL U_g1768 (.A(G947_1353_gat), .Y(G947_1353_ngat) );
INVXL U_g1769 (.A(G948_1319_gat), .Y(G948_1319_ngat) );
INVXL U_g1770 (.A(G955_1351_gat), .Y(G955_1351_ngat) );
INVXL U_g1771 (.A(G956_1321_gat), .Y(G956_1321_ngat) );
INVXL U_g1772 (.A(G1165_1356_gat), .Y(G1165_1356_ngat) );
INVXL U_g1773 (.A(G1166_1325_gat), .Y(G1166_1325_ngat) );
INVXL U_g1774 (.A(G1173_1354_gat), .Y(G1173_1354_ngat) );
INVXL U_g1775 (.A(G1174_1327_gat), .Y(G1174_1327_ngat) );
INVXL U_g1776 (.A(G641_1365_gat), .Y(G641_1365_ngat) );
INVXL U_g1777 (.A(G642_1345_gat), .Y(G642_1345_ngat) );
INVXL U_g1778 (.A(G648_1366_gat), .Y(G648_1366_ngat) );
INVXL U_g1779 (.A(G649_1346_gat), .Y(G649_1346_ngat) );
INVXL U_g1780 (.A(G976_1373_gat), .Y(G976_1373_ngat) );
INVXL U_g1781 (.A(G969_1359_gat), .Y(G969_1359_ngat) );
INVXL U_g1782 (.A(G1193_1374_gat), .Y(G1193_1374_ngat) );
INVXL U_g1783 (.A(G1186_1360_gat), .Y(G1186_1360_ngat) );
INVXL U_g1784 (.A(G329_1414_gat), .Y(G329_1414_ngat) );
INVXL U_g1785 (.A(G991_1411_gat), .Y(G991_1411_ngat) );

endmodule
