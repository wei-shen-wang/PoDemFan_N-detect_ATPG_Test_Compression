module C6288 ( G1GAT_0_gat, G18GAT_1_gat, G35GAT_2_gat, G52GAT_3_gat, G69GAT_4_gat, G86GAT_5_gat, G103GAT_6_gat, G120GAT_7_gat, G137GAT_8_gat, G154GAT_9_gat, G171GAT_10_gat, G188GAT_11_gat, G205GAT_12_gat, G222GAT_13_gat, G239GAT_14_gat, G256GAT_15_gat, G273GAT_16_gat, G290GAT_17_gat, G307GAT_18_gat, G324GAT_19_gat, G341GAT_20_gat, G358GAT_21_gat, G375GAT_22_gat, G392GAT_23_gat, G409GAT_24_gat, G426GAT_25_gat, G443GAT_26_gat, G460GAT_27_gat, G477GAT_28_gat, G494GAT_29_gat, G511GAT_30_gat, G528GAT_31_gat, G545GAT_287_gat, G1581GAT_423_gat, G1901GAT_561_gat, G2223GAT_700_gat, G2548GAT_840_gat, G2877GAT_983_gat, G3211GAT_1128_gat, G3552GAT_1275_gat, G3895GAT_1423_gat, G4241GAT_1572_gat, G4591GAT_1722_gat, G4946GAT_1876_gat, G5308GAT_2031_gat, G5672GAT_2187_gat, G5971GAT_2309_gat, G6123GAT_2368_gat, G6150GAT_2378_gat, G6160GAT_2383_gat, G6170GAT_2388_gat, G6180GAT_2393_gat, G6190GAT_2398_gat, G6200GAT_2403_gat, G6210GAT_2408_gat, G6220GAT_2413_gat, G6230GAT_2418_gat, G6240GAT_2423_gat, G6250GAT_2428_gat, G6260GAT_2433_gat, G6270GAT_2438_gat, G6280GAT_2443_gat, G6287GAT_2444_gat, G6288GAT_2447_gat);

input G1GAT_0_gat;
input G18GAT_1_gat;
input G35GAT_2_gat;
input G52GAT_3_gat;
input G69GAT_4_gat;
input G86GAT_5_gat;
input G103GAT_6_gat;
input G120GAT_7_gat;
input G137GAT_8_gat;
input G154GAT_9_gat;
input G171GAT_10_gat;
input G188GAT_11_gat;
input G205GAT_12_gat;
input G222GAT_13_gat;
input G239GAT_14_gat;
input G256GAT_15_gat;
input G273GAT_16_gat;
input G290GAT_17_gat;
input G307GAT_18_gat;
input G324GAT_19_gat;
input G341GAT_20_gat;
input G358GAT_21_gat;
input G375GAT_22_gat;
input G392GAT_23_gat;
input G409GAT_24_gat;
input G426GAT_25_gat;
input G443GAT_26_gat;
input G460GAT_27_gat;
input G477GAT_28_gat;
input G494GAT_29_gat;
input G511GAT_30_gat;
input G528GAT_31_gat;

output G545GAT_287_gat;
output G1581GAT_423_gat;
output G1901GAT_561_gat;
output G2223GAT_700_gat;
output G2548GAT_840_gat;
output G2877GAT_983_gat;
output G3211GAT_1128_gat;
output G3552GAT_1275_gat;
output G3895GAT_1423_gat;
output G4241GAT_1572_gat;
output G4591GAT_1722_gat;
output G4946GAT_1876_gat;
output G5308GAT_2031_gat;
output G5672GAT_2187_gat;
output G5971GAT_2309_gat;
output G6123GAT_2368_gat;
output G6150GAT_2378_gat;
output G6160GAT_2383_gat;
output G6170GAT_2388_gat;
output G6180GAT_2393_gat;
output G6190GAT_2398_gat;
output G6200GAT_2403_gat;
output G6210GAT_2408_gat;
output G6220GAT_2413_gat;
output G6230GAT_2418_gat;
output G6240GAT_2423_gat;
output G6250GAT_2428_gat;
output G6260GAT_2433_gat;
output G6270GAT_2438_gat;
output G6280GAT_2443_gat;
output G6287GAT_2444_gat;
output G6288GAT_2447_gat;

AND2XL U_g1 (.A(G528GAT_31_gat), .B(G256GAT_15_gat), .Y(G1308GAT_32_gat) );
AND2XL U_g2 (.A(G511GAT_30_gat), .B(G256GAT_15_gat), .Y(G1305GAT_33_gat) );
AND2XL U_g3 (.A(G494GAT_29_gat), .B(G256GAT_15_gat), .Y(G1302GAT_34_gat) );
AND2XL U_g4 (.A(G477GAT_28_gat), .B(G256GAT_15_gat), .Y(G1299GAT_35_gat) );
AND2XL U_g5 (.A(G460GAT_27_gat), .B(G256GAT_15_gat), .Y(G1296GAT_36_gat) );
AND2XL U_g6 (.A(G443GAT_26_gat), .B(G256GAT_15_gat), .Y(G1293GAT_37_gat) );
AND2XL U_g7 (.A(G426GAT_25_gat), .B(G256GAT_15_gat), .Y(G1290GAT_38_gat) );
AND2XL U_g8 (.A(G409GAT_24_gat), .B(G256GAT_15_gat), .Y(G1287GAT_39_gat) );
AND2XL U_g9 (.A(G392GAT_23_gat), .B(G256GAT_15_gat), .Y(G1284GAT_40_gat) );
AND2XL U_g10 (.A(G375GAT_22_gat), .B(G256GAT_15_gat), .Y(G1281GAT_41_gat) );
AND2XL U_g11 (.A(G358GAT_21_gat), .B(G256GAT_15_gat), .Y(G1278GAT_42_gat) );
AND2XL U_g12 (.A(G341GAT_20_gat), .B(G256GAT_15_gat), .Y(G1275GAT_43_gat) );
AND2XL U_g13 (.A(G324GAT_19_gat), .B(G256GAT_15_gat), .Y(G1272GAT_44_gat) );
AND2XL U_g14 (.A(G307GAT_18_gat), .B(G256GAT_15_gat), .Y(G1269GAT_45_gat) );
AND2XL U_g15 (.A(G290GAT_17_gat), .B(G256GAT_15_gat), .Y(G1266GAT_46_gat) );
AND2XL U_g16 (.A(G273GAT_16_gat), .B(G256GAT_15_gat), .Y(G1263GAT_47_gat) );
AND2XL U_g17 (.A(G528GAT_31_gat), .B(G239GAT_14_gat), .Y(G1260GAT_48_gat) );
AND2XL U_g18 (.A(G511GAT_30_gat), .B(G239GAT_14_gat), .Y(G1257GAT_49_gat) );
AND2XL U_g19 (.A(G494GAT_29_gat), .B(G239GAT_14_gat), .Y(G1254GAT_50_gat) );
AND2XL U_g20 (.A(G477GAT_28_gat), .B(G239GAT_14_gat), .Y(G1251GAT_51_gat) );
AND2XL U_g21 (.A(G460GAT_27_gat), .B(G239GAT_14_gat), .Y(G1248GAT_52_gat) );
AND2XL U_g22 (.A(G443GAT_26_gat), .B(G239GAT_14_gat), .Y(G1245GAT_53_gat) );
AND2XL U_g23 (.A(G426GAT_25_gat), .B(G239GAT_14_gat), .Y(G1242GAT_54_gat) );
AND2XL U_g24 (.A(G409GAT_24_gat), .B(G239GAT_14_gat), .Y(G1239GAT_55_gat) );
AND2XL U_g25 (.A(G392GAT_23_gat), .B(G239GAT_14_gat), .Y(G1236GAT_56_gat) );
AND2XL U_g26 (.A(G375GAT_22_gat), .B(G239GAT_14_gat), .Y(G1233GAT_57_gat) );
AND2XL U_g27 (.A(G358GAT_21_gat), .B(G239GAT_14_gat), .Y(G1230GAT_58_gat) );
AND2XL U_g28 (.A(G341GAT_20_gat), .B(G239GAT_14_gat), .Y(G1227GAT_59_gat) );
AND2XL U_g29 (.A(G324GAT_19_gat), .B(G239GAT_14_gat), .Y(G1224GAT_60_gat) );
AND2XL U_g30 (.A(G307GAT_18_gat), .B(G239GAT_14_gat), .Y(G1221GAT_61_gat) );
AND2XL U_g31 (.A(G290GAT_17_gat), .B(G239GAT_14_gat), .Y(G1218GAT_62_gat) );
AND2XL U_g32 (.A(G273GAT_16_gat), .B(G239GAT_14_gat), .Y(G1215GAT_63_gat) );
AND2XL U_g33 (.A(G528GAT_31_gat), .B(G222GAT_13_gat), .Y(G1212GAT_64_gat) );
AND2XL U_g34 (.A(G511GAT_30_gat), .B(G222GAT_13_gat), .Y(G1209GAT_65_gat) );
AND2XL U_g35 (.A(G494GAT_29_gat), .B(G222GAT_13_gat), .Y(G1206GAT_66_gat) );
AND2XL U_g36 (.A(G477GAT_28_gat), .B(G222GAT_13_gat), .Y(G1203GAT_67_gat) );
AND2XL U_g37 (.A(G460GAT_27_gat), .B(G222GAT_13_gat), .Y(G1200GAT_68_gat) );
AND2XL U_g38 (.A(G443GAT_26_gat), .B(G222GAT_13_gat), .Y(G1197GAT_69_gat) );
AND2XL U_g39 (.A(G426GAT_25_gat), .B(G222GAT_13_gat), .Y(G1194GAT_70_gat) );
AND2XL U_g40 (.A(G409GAT_24_gat), .B(G222GAT_13_gat), .Y(G1191GAT_71_gat) );
AND2XL U_g41 (.A(G392GAT_23_gat), .B(G222GAT_13_gat), .Y(G1188GAT_72_gat) );
AND2XL U_g42 (.A(G375GAT_22_gat), .B(G222GAT_13_gat), .Y(G1185GAT_73_gat) );
AND2XL U_g43 (.A(G358GAT_21_gat), .B(G222GAT_13_gat), .Y(G1182GAT_74_gat) );
AND2XL U_g44 (.A(G341GAT_20_gat), .B(G222GAT_13_gat), .Y(G1179GAT_75_gat) );
AND2XL U_g45 (.A(G324GAT_19_gat), .B(G222GAT_13_gat), .Y(G1176GAT_76_gat) );
AND2XL U_g46 (.A(G307GAT_18_gat), .B(G222GAT_13_gat), .Y(G1173GAT_77_gat) );
AND2XL U_g47 (.A(G290GAT_17_gat), .B(G222GAT_13_gat), .Y(G1170GAT_78_gat) );
AND2XL U_g48 (.A(G273GAT_16_gat), .B(G222GAT_13_gat), .Y(G1167GAT_79_gat) );
AND2XL U_g49 (.A(G528GAT_31_gat), .B(G205GAT_12_gat), .Y(G1164GAT_80_gat) );
AND2XL U_g50 (.A(G511GAT_30_gat), .B(G205GAT_12_gat), .Y(G1161GAT_81_gat) );
AND2XL U_g51 (.A(G494GAT_29_gat), .B(G205GAT_12_gat), .Y(G1158GAT_82_gat) );
AND2XL U_g52 (.A(G477GAT_28_gat), .B(G205GAT_12_gat), .Y(G1155GAT_83_gat) );
AND2XL U_g53 (.A(G460GAT_27_gat), .B(G205GAT_12_gat), .Y(G1152GAT_84_gat) );
AND2XL U_g54 (.A(G443GAT_26_gat), .B(G205GAT_12_gat), .Y(G1149GAT_85_gat) );
AND2XL U_g55 (.A(G426GAT_25_gat), .B(G205GAT_12_gat), .Y(G1146GAT_86_gat) );
AND2XL U_g56 (.A(G409GAT_24_gat), .B(G205GAT_12_gat), .Y(G1143GAT_87_gat) );
AND2XL U_g57 (.A(G392GAT_23_gat), .B(G205GAT_12_gat), .Y(G1140GAT_88_gat) );
AND2XL U_g58 (.A(G375GAT_22_gat), .B(G205GAT_12_gat), .Y(G1137GAT_89_gat) );
AND2XL U_g59 (.A(G358GAT_21_gat), .B(G205GAT_12_gat), .Y(G1134GAT_90_gat) );
AND2XL U_g60 (.A(G341GAT_20_gat), .B(G205GAT_12_gat), .Y(G1131GAT_91_gat) );
AND2XL U_g61 (.A(G324GAT_19_gat), .B(G205GAT_12_gat), .Y(G1128GAT_92_gat) );
AND2XL U_g62 (.A(G307GAT_18_gat), .B(G205GAT_12_gat), .Y(G1125GAT_93_gat) );
AND2XL U_g63 (.A(G290GAT_17_gat), .B(G205GAT_12_gat), .Y(G1122GAT_94_gat) );
AND2XL U_g64 (.A(G273GAT_16_gat), .B(G205GAT_12_gat), .Y(G1119GAT_95_gat) );
AND2XL U_g65 (.A(G528GAT_31_gat), .B(G188GAT_11_gat), .Y(G1116GAT_96_gat) );
AND2XL U_g66 (.A(G511GAT_30_gat), .B(G188GAT_11_gat), .Y(G1113GAT_97_gat) );
AND2XL U_g67 (.A(G494GAT_29_gat), .B(G188GAT_11_gat), .Y(G1110GAT_98_gat) );
AND2XL U_g68 (.A(G477GAT_28_gat), .B(G188GAT_11_gat), .Y(G1107GAT_99_gat) );
AND2XL U_g69 (.A(G460GAT_27_gat), .B(G188GAT_11_gat), .Y(G1104GAT_100_gat) );
AND2XL U_g70 (.A(G443GAT_26_gat), .B(G188GAT_11_gat), .Y(G1101GAT_101_gat) );
AND2XL U_g71 (.A(G426GAT_25_gat), .B(G188GAT_11_gat), .Y(G1098GAT_102_gat) );
AND2XL U_g72 (.A(G409GAT_24_gat), .B(G188GAT_11_gat), .Y(G1095GAT_103_gat) );
AND2XL U_g73 (.A(G392GAT_23_gat), .B(G188GAT_11_gat), .Y(G1092GAT_104_gat) );
AND2XL U_g74 (.A(G375GAT_22_gat), .B(G188GAT_11_gat), .Y(G1089GAT_105_gat) );
AND2XL U_g75 (.A(G358GAT_21_gat), .B(G188GAT_11_gat), .Y(G1086GAT_106_gat) );
AND2XL U_g76 (.A(G341GAT_20_gat), .B(G188GAT_11_gat), .Y(G1083GAT_107_gat) );
AND2XL U_g77 (.A(G324GAT_19_gat), .B(G188GAT_11_gat), .Y(G1080GAT_108_gat) );
AND2XL U_g78 (.A(G307GAT_18_gat), .B(G188GAT_11_gat), .Y(G1077GAT_109_gat) );
AND2XL U_g79 (.A(G290GAT_17_gat), .B(G188GAT_11_gat), .Y(G1074GAT_110_gat) );
AND2XL U_g80 (.A(G273GAT_16_gat), .B(G188GAT_11_gat), .Y(G1071GAT_111_gat) );
AND2XL U_g81 (.A(G528GAT_31_gat), .B(G171GAT_10_gat), .Y(G1068GAT_112_gat) );
AND2XL U_g82 (.A(G511GAT_30_gat), .B(G171GAT_10_gat), .Y(G1065GAT_113_gat) );
AND2XL U_g83 (.A(G494GAT_29_gat), .B(G171GAT_10_gat), .Y(G1062GAT_114_gat) );
AND2XL U_g84 (.A(G477GAT_28_gat), .B(G171GAT_10_gat), .Y(G1059GAT_115_gat) );
AND2XL U_g85 (.A(G460GAT_27_gat), .B(G171GAT_10_gat), .Y(G1056GAT_116_gat) );
AND2XL U_g86 (.A(G443GAT_26_gat), .B(G171GAT_10_gat), .Y(G1053GAT_117_gat) );
AND2XL U_g87 (.A(G426GAT_25_gat), .B(G171GAT_10_gat), .Y(G1050GAT_118_gat) );
AND2XL U_g88 (.A(G409GAT_24_gat), .B(G171GAT_10_gat), .Y(G1047GAT_119_gat) );
AND2XL U_g89 (.A(G392GAT_23_gat), .B(G171GAT_10_gat), .Y(G1044GAT_120_gat) );
AND2XL U_g90 (.A(G375GAT_22_gat), .B(G171GAT_10_gat), .Y(G1041GAT_121_gat) );
AND2XL U_g91 (.A(G358GAT_21_gat), .B(G171GAT_10_gat), .Y(G1038GAT_122_gat) );
AND2XL U_g92 (.A(G341GAT_20_gat), .B(G171GAT_10_gat), .Y(G1035GAT_123_gat) );
AND2XL U_g93 (.A(G324GAT_19_gat), .B(G171GAT_10_gat), .Y(G1032GAT_124_gat) );
AND2XL U_g94 (.A(G307GAT_18_gat), .B(G171GAT_10_gat), .Y(G1029GAT_125_gat) );
AND2XL U_g95 (.A(G290GAT_17_gat), .B(G171GAT_10_gat), .Y(G1026GAT_126_gat) );
AND2XL U_g96 (.A(G273GAT_16_gat), .B(G171GAT_10_gat), .Y(G1023GAT_127_gat) );
AND2XL U_g97 (.A(G528GAT_31_gat), .B(G154GAT_9_gat), .Y(G1020GAT_128_gat) );
AND2XL U_g98 (.A(G511GAT_30_gat), .B(G154GAT_9_gat), .Y(G1017GAT_129_gat) );
AND2XL U_g99 (.A(G494GAT_29_gat), .B(G154GAT_9_gat), .Y(G1014GAT_130_gat) );
AND2XL U_g100 (.A(G477GAT_28_gat), .B(G154GAT_9_gat), .Y(G1011GAT_131_gat) );
AND2XL U_g101 (.A(G460GAT_27_gat), .B(G154GAT_9_gat), .Y(G1008GAT_132_gat) );
AND2XL U_g102 (.A(G443GAT_26_gat), .B(G154GAT_9_gat), .Y(G1005GAT_133_gat) );
AND2XL U_g103 (.A(G426GAT_25_gat), .B(G154GAT_9_gat), .Y(G1002GAT_134_gat) );
AND2XL U_g104 (.A(G409GAT_24_gat), .B(G154GAT_9_gat), .Y(G999GAT_135_gat) );
AND2XL U_g105 (.A(G392GAT_23_gat), .B(G154GAT_9_gat), .Y(G996GAT_136_gat) );
AND2XL U_g106 (.A(G375GAT_22_gat), .B(G154GAT_9_gat), .Y(G993GAT_137_gat) );
AND2XL U_g107 (.A(G358GAT_21_gat), .B(G154GAT_9_gat), .Y(G990GAT_138_gat) );
AND2XL U_g108 (.A(G341GAT_20_gat), .B(G154GAT_9_gat), .Y(G987GAT_139_gat) );
AND2XL U_g109 (.A(G324GAT_19_gat), .B(G154GAT_9_gat), .Y(G984GAT_140_gat) );
AND2XL U_g110 (.A(G307GAT_18_gat), .B(G154GAT_9_gat), .Y(G981GAT_141_gat) );
AND2XL U_g111 (.A(G290GAT_17_gat), .B(G154GAT_9_gat), .Y(G978GAT_142_gat) );
AND2XL U_g112 (.A(G273GAT_16_gat), .B(G154GAT_9_gat), .Y(G975GAT_143_gat) );
AND2XL U_g113 (.A(G528GAT_31_gat), .B(G137GAT_8_gat), .Y(G972GAT_144_gat) );
AND2XL U_g114 (.A(G511GAT_30_gat), .B(G137GAT_8_gat), .Y(G969GAT_145_gat) );
AND2XL U_g115 (.A(G494GAT_29_gat), .B(G137GAT_8_gat), .Y(G966GAT_146_gat) );
AND2XL U_g116 (.A(G477GAT_28_gat), .B(G137GAT_8_gat), .Y(G963GAT_147_gat) );
AND2XL U_g117 (.A(G460GAT_27_gat), .B(G137GAT_8_gat), .Y(G960GAT_148_gat) );
AND2XL U_g118 (.A(G443GAT_26_gat), .B(G137GAT_8_gat), .Y(G957GAT_149_gat) );
AND2XL U_g119 (.A(G426GAT_25_gat), .B(G137GAT_8_gat), .Y(G954GAT_150_gat) );
AND2XL U_g120 (.A(G409GAT_24_gat), .B(G137GAT_8_gat), .Y(G951GAT_151_gat) );
AND2XL U_g121 (.A(G392GAT_23_gat), .B(G137GAT_8_gat), .Y(G948GAT_152_gat) );
AND2XL U_g122 (.A(G375GAT_22_gat), .B(G137GAT_8_gat), .Y(G945GAT_153_gat) );
AND2XL U_g123 (.A(G358GAT_21_gat), .B(G137GAT_8_gat), .Y(G942GAT_154_gat) );
AND2XL U_g124 (.A(G341GAT_20_gat), .B(G137GAT_8_gat), .Y(G939GAT_155_gat) );
AND2XL U_g125 (.A(G324GAT_19_gat), .B(G137GAT_8_gat), .Y(G936GAT_156_gat) );
AND2XL U_g126 (.A(G307GAT_18_gat), .B(G137GAT_8_gat), .Y(G933GAT_157_gat) );
AND2XL U_g127 (.A(G290GAT_17_gat), .B(G137GAT_8_gat), .Y(G930GAT_158_gat) );
AND2XL U_g128 (.A(G273GAT_16_gat), .B(G137GAT_8_gat), .Y(G927GAT_159_gat) );
AND2XL U_g129 (.A(G528GAT_31_gat), .B(G120GAT_7_gat), .Y(G924GAT_160_gat) );
AND2XL U_g130 (.A(G511GAT_30_gat), .B(G120GAT_7_gat), .Y(G921GAT_161_gat) );
AND2XL U_g131 (.A(G494GAT_29_gat), .B(G120GAT_7_gat), .Y(G918GAT_162_gat) );
AND2XL U_g132 (.A(G477GAT_28_gat), .B(G120GAT_7_gat), .Y(G915GAT_163_gat) );
AND2XL U_g133 (.A(G460GAT_27_gat), .B(G120GAT_7_gat), .Y(G912GAT_164_gat) );
AND2XL U_g134 (.A(G443GAT_26_gat), .B(G120GAT_7_gat), .Y(G909GAT_165_gat) );
AND2XL U_g135 (.A(G426GAT_25_gat), .B(G120GAT_7_gat), .Y(G906GAT_166_gat) );
AND2XL U_g136 (.A(G409GAT_24_gat), .B(G120GAT_7_gat), .Y(G903GAT_167_gat) );
AND2XL U_g137 (.A(G392GAT_23_gat), .B(G120GAT_7_gat), .Y(G900GAT_168_gat) );
AND2XL U_g138 (.A(G375GAT_22_gat), .B(G120GAT_7_gat), .Y(G897GAT_169_gat) );
AND2XL U_g139 (.A(G358GAT_21_gat), .B(G120GAT_7_gat), .Y(G894GAT_170_gat) );
AND2XL U_g140 (.A(G341GAT_20_gat), .B(G120GAT_7_gat), .Y(G891GAT_171_gat) );
AND2XL U_g141 (.A(G324GAT_19_gat), .B(G120GAT_7_gat), .Y(G888GAT_172_gat) );
AND2XL U_g142 (.A(G307GAT_18_gat), .B(G120GAT_7_gat), .Y(G885GAT_173_gat) );
AND2XL U_g143 (.A(G290GAT_17_gat), .B(G120GAT_7_gat), .Y(G882GAT_174_gat) );
AND2XL U_g144 (.A(G273GAT_16_gat), .B(G120GAT_7_gat), .Y(G879GAT_175_gat) );
AND2XL U_g145 (.A(G528GAT_31_gat), .B(G103GAT_6_gat), .Y(G876GAT_176_gat) );
AND2XL U_g146 (.A(G511GAT_30_gat), .B(G103GAT_6_gat), .Y(G873GAT_177_gat) );
AND2XL U_g147 (.A(G494GAT_29_gat), .B(G103GAT_6_gat), .Y(G870GAT_178_gat) );
AND2XL U_g148 (.A(G477GAT_28_gat), .B(G103GAT_6_gat), .Y(G867GAT_179_gat) );
AND2XL U_g149 (.A(G460GAT_27_gat), .B(G103GAT_6_gat), .Y(G864GAT_180_gat) );
AND2XL U_g150 (.A(G443GAT_26_gat), .B(G103GAT_6_gat), .Y(G861GAT_181_gat) );
AND2XL U_g151 (.A(G426GAT_25_gat), .B(G103GAT_6_gat), .Y(G858GAT_182_gat) );
AND2XL U_g152 (.A(G409GAT_24_gat), .B(G103GAT_6_gat), .Y(G855GAT_183_gat) );
AND2XL U_g153 (.A(G392GAT_23_gat), .B(G103GAT_6_gat), .Y(G852GAT_184_gat) );
AND2XL U_g154 (.A(G375GAT_22_gat), .B(G103GAT_6_gat), .Y(G849GAT_185_gat) );
AND2XL U_g155 (.A(G358GAT_21_gat), .B(G103GAT_6_gat), .Y(G846GAT_186_gat) );
AND2XL U_g156 (.A(G341GAT_20_gat), .B(G103GAT_6_gat), .Y(G843GAT_187_gat) );
AND2XL U_g157 (.A(G324GAT_19_gat), .B(G103GAT_6_gat), .Y(G840GAT_188_gat) );
AND2XL U_g158 (.A(G307GAT_18_gat), .B(G103GAT_6_gat), .Y(G837GAT_189_gat) );
AND2XL U_g159 (.A(G290GAT_17_gat), .B(G103GAT_6_gat), .Y(G834GAT_190_gat) );
AND2XL U_g160 (.A(G273GAT_16_gat), .B(G103GAT_6_gat), .Y(G831GAT_191_gat) );
AND2XL U_g161 (.A(G528GAT_31_gat), .B(G86GAT_5_gat), .Y(G828GAT_192_gat) );
AND2XL U_g162 (.A(G511GAT_30_gat), .B(G86GAT_5_gat), .Y(G825GAT_193_gat) );
AND2XL U_g163 (.A(G494GAT_29_gat), .B(G86GAT_5_gat), .Y(G822GAT_194_gat) );
AND2XL U_g164 (.A(G477GAT_28_gat), .B(G86GAT_5_gat), .Y(G819GAT_195_gat) );
AND2XL U_g165 (.A(G460GAT_27_gat), .B(G86GAT_5_gat), .Y(G816GAT_196_gat) );
AND2XL U_g166 (.A(G443GAT_26_gat), .B(G86GAT_5_gat), .Y(G813GAT_197_gat) );
AND2XL U_g167 (.A(G426GAT_25_gat), .B(G86GAT_5_gat), .Y(G810GAT_198_gat) );
AND2XL U_g168 (.A(G409GAT_24_gat), .B(G86GAT_5_gat), .Y(G807GAT_199_gat) );
AND2XL U_g169 (.A(G392GAT_23_gat), .B(G86GAT_5_gat), .Y(G804GAT_200_gat) );
AND2XL U_g170 (.A(G375GAT_22_gat), .B(G86GAT_5_gat), .Y(G801GAT_201_gat) );
AND2XL U_g171 (.A(G358GAT_21_gat), .B(G86GAT_5_gat), .Y(G798GAT_202_gat) );
AND2XL U_g172 (.A(G341GAT_20_gat), .B(G86GAT_5_gat), .Y(G795GAT_203_gat) );
AND2XL U_g173 (.A(G324GAT_19_gat), .B(G86GAT_5_gat), .Y(G792GAT_204_gat) );
AND2XL U_g174 (.A(G307GAT_18_gat), .B(G86GAT_5_gat), .Y(G789GAT_205_gat) );
AND2XL U_g175 (.A(G290GAT_17_gat), .B(G86GAT_5_gat), .Y(G786GAT_206_gat) );
AND2XL U_g176 (.A(G273GAT_16_gat), .B(G86GAT_5_gat), .Y(G783GAT_207_gat) );
AND2XL U_g177 (.A(G528GAT_31_gat), .B(G69GAT_4_gat), .Y(G780GAT_208_gat) );
AND2XL U_g178 (.A(G511GAT_30_gat), .B(G69GAT_4_gat), .Y(G777GAT_209_gat) );
AND2XL U_g179 (.A(G494GAT_29_gat), .B(G69GAT_4_gat), .Y(G774GAT_210_gat) );
AND2XL U_g180 (.A(G477GAT_28_gat), .B(G69GAT_4_gat), .Y(G771GAT_211_gat) );
AND2XL U_g181 (.A(G460GAT_27_gat), .B(G69GAT_4_gat), .Y(G768GAT_212_gat) );
AND2XL U_g182 (.A(G443GAT_26_gat), .B(G69GAT_4_gat), .Y(G765GAT_213_gat) );
AND2XL U_g183 (.A(G426GAT_25_gat), .B(G69GAT_4_gat), .Y(G762GAT_214_gat) );
AND2XL U_g184 (.A(G409GAT_24_gat), .B(G69GAT_4_gat), .Y(G759GAT_215_gat) );
AND2XL U_g185 (.A(G392GAT_23_gat), .B(G69GAT_4_gat), .Y(G756GAT_216_gat) );
AND2XL U_g186 (.A(G375GAT_22_gat), .B(G69GAT_4_gat), .Y(G753GAT_217_gat) );
AND2XL U_g187 (.A(G358GAT_21_gat), .B(G69GAT_4_gat), .Y(G750GAT_218_gat) );
AND2XL U_g188 (.A(G341GAT_20_gat), .B(G69GAT_4_gat), .Y(G747GAT_219_gat) );
AND2XL U_g189 (.A(G324GAT_19_gat), .B(G69GAT_4_gat), .Y(G744GAT_220_gat) );
AND2XL U_g190 (.A(G307GAT_18_gat), .B(G69GAT_4_gat), .Y(G741GAT_221_gat) );
AND2XL U_g191 (.A(G290GAT_17_gat), .B(G69GAT_4_gat), .Y(G738GAT_222_gat) );
AND2XL U_g192 (.A(G273GAT_16_gat), .B(G69GAT_4_gat), .Y(G735GAT_223_gat) );
AND2XL U_g193 (.A(G528GAT_31_gat), .B(G52GAT_3_gat), .Y(G732GAT_224_gat) );
AND2XL U_g194 (.A(G511GAT_30_gat), .B(G52GAT_3_gat), .Y(G729GAT_225_gat) );
AND2XL U_g195 (.A(G494GAT_29_gat), .B(G52GAT_3_gat), .Y(G726GAT_226_gat) );
AND2XL U_g196 (.A(G477GAT_28_gat), .B(G52GAT_3_gat), .Y(G723GAT_227_gat) );
AND2XL U_g197 (.A(G460GAT_27_gat), .B(G52GAT_3_gat), .Y(G720GAT_228_gat) );
AND2XL U_g198 (.A(G443GAT_26_gat), .B(G52GAT_3_gat), .Y(G717GAT_229_gat) );
AND2XL U_g199 (.A(G426GAT_25_gat), .B(G52GAT_3_gat), .Y(G714GAT_230_gat) );
AND2XL U_g200 (.A(G409GAT_24_gat), .B(G52GAT_3_gat), .Y(G711GAT_231_gat) );
AND2XL U_g201 (.A(G392GAT_23_gat), .B(G52GAT_3_gat), .Y(G708GAT_232_gat) );
AND2XL U_g202 (.A(G375GAT_22_gat), .B(G52GAT_3_gat), .Y(G705GAT_233_gat) );
AND2XL U_g203 (.A(G358GAT_21_gat), .B(G52GAT_3_gat), .Y(G702GAT_234_gat) );
AND2XL U_g204 (.A(G341GAT_20_gat), .B(G52GAT_3_gat), .Y(G699GAT_235_gat) );
AND2XL U_g205 (.A(G324GAT_19_gat), .B(G52GAT_3_gat), .Y(G696GAT_236_gat) );
AND2XL U_g206 (.A(G307GAT_18_gat), .B(G52GAT_3_gat), .Y(G693GAT_237_gat) );
AND2XL U_g207 (.A(G290GAT_17_gat), .B(G52GAT_3_gat), .Y(G690GAT_238_gat) );
AND2XL U_g208 (.A(G273GAT_16_gat), .B(G52GAT_3_gat), .Y(G687GAT_239_gat) );
AND2XL U_g209 (.A(G528GAT_31_gat), .B(G35GAT_2_gat), .Y(G684GAT_240_gat) );
AND2XL U_g210 (.A(G511GAT_30_gat), .B(G35GAT_2_gat), .Y(G681GAT_241_gat) );
AND2XL U_g211 (.A(G494GAT_29_gat), .B(G35GAT_2_gat), .Y(G678GAT_242_gat) );
AND2XL U_g212 (.A(G477GAT_28_gat), .B(G35GAT_2_gat), .Y(G675GAT_243_gat) );
AND2XL U_g213 (.A(G460GAT_27_gat), .B(G35GAT_2_gat), .Y(G672GAT_244_gat) );
AND2XL U_g214 (.A(G443GAT_26_gat), .B(G35GAT_2_gat), .Y(G669GAT_245_gat) );
AND2XL U_g215 (.A(G426GAT_25_gat), .B(G35GAT_2_gat), .Y(G666GAT_246_gat) );
AND2XL U_g216 (.A(G409GAT_24_gat), .B(G35GAT_2_gat), .Y(G663GAT_247_gat) );
AND2XL U_g217 (.A(G392GAT_23_gat), .B(G35GAT_2_gat), .Y(G660GAT_248_gat) );
AND2XL U_g218 (.A(G375GAT_22_gat), .B(G35GAT_2_gat), .Y(G657GAT_249_gat) );
AND2XL U_g219 (.A(G358GAT_21_gat), .B(G35GAT_2_gat), .Y(G654GAT_250_gat) );
AND2XL U_g220 (.A(G341GAT_20_gat), .B(G35GAT_2_gat), .Y(G651GAT_251_gat) );
AND2XL U_g221 (.A(G324GAT_19_gat), .B(G35GAT_2_gat), .Y(G648GAT_252_gat) );
AND2XL U_g222 (.A(G307GAT_18_gat), .B(G35GAT_2_gat), .Y(G645GAT_253_gat) );
AND2XL U_g223 (.A(G290GAT_17_gat), .B(G35GAT_2_gat), .Y(G642GAT_254_gat) );
AND2XL U_g224 (.A(G273GAT_16_gat), .B(G35GAT_2_gat), .Y(G639GAT_255_gat) );
AND2XL U_g225 (.A(G528GAT_31_gat), .B(G18GAT_1_gat), .Y(G636GAT_256_gat) );
AND2XL U_g226 (.A(G511GAT_30_gat), .B(G18GAT_1_gat), .Y(G633GAT_257_gat) );
AND2XL U_g227 (.A(G494GAT_29_gat), .B(G18GAT_1_gat), .Y(G630GAT_258_gat) );
AND2XL U_g228 (.A(G477GAT_28_gat), .B(G18GAT_1_gat), .Y(G627GAT_259_gat) );
AND2XL U_g229 (.A(G460GAT_27_gat), .B(G18GAT_1_gat), .Y(G624GAT_260_gat) );
AND2XL U_g230 (.A(G443GAT_26_gat), .B(G18GAT_1_gat), .Y(G621GAT_261_gat) );
AND2XL U_g231 (.A(G426GAT_25_gat), .B(G18GAT_1_gat), .Y(G618GAT_262_gat) );
AND2XL U_g232 (.A(G409GAT_24_gat), .B(G18GAT_1_gat), .Y(G615GAT_263_gat) );
AND2XL U_g233 (.A(G392GAT_23_gat), .B(G18GAT_1_gat), .Y(G612GAT_264_gat) );
AND2XL U_g234 (.A(G375GAT_22_gat), .B(G18GAT_1_gat), .Y(G609GAT_265_gat) );
AND2XL U_g235 (.A(G358GAT_21_gat), .B(G18GAT_1_gat), .Y(G606GAT_266_gat) );
AND2XL U_g236 (.A(G341GAT_20_gat), .B(G18GAT_1_gat), .Y(G603GAT_267_gat) );
AND2XL U_g237 (.A(G324GAT_19_gat), .B(G18GAT_1_gat), .Y(G600GAT_268_gat) );
AND2XL U_g238 (.A(G307GAT_18_gat), .B(G18GAT_1_gat), .Y(G597GAT_269_gat) );
AND2XL U_g239 (.A(G290GAT_17_gat), .B(G18GAT_1_gat), .Y(G594GAT_270_gat) );
AND2XL U_g240 (.A(G273GAT_16_gat), .B(G18GAT_1_gat), .Y(G591GAT_271_gat) );
AND2XL U_g241 (.A(G528GAT_31_gat), .B(G1GAT_0_gat), .Y(G588GAT_272_gat) );
AND2XL U_g242 (.A(G511GAT_30_gat), .B(G1GAT_0_gat), .Y(G585GAT_273_gat) );
AND2XL U_g243 (.A(G494GAT_29_gat), .B(G1GAT_0_gat), .Y(G582GAT_274_gat) );
AND2XL U_g244 (.A(G477GAT_28_gat), .B(G1GAT_0_gat), .Y(G579GAT_275_gat) );
AND2XL U_g245 (.A(G460GAT_27_gat), .B(G1GAT_0_gat), .Y(G576GAT_276_gat) );
AND2XL U_g246 (.A(G443GAT_26_gat), .B(G1GAT_0_gat), .Y(G573GAT_277_gat) );
AND2XL U_g247 (.A(G426GAT_25_gat), .B(G1GAT_0_gat), .Y(G570GAT_278_gat) );
AND2XL U_g248 (.A(G409GAT_24_gat), .B(G1GAT_0_gat), .Y(G567GAT_279_gat) );
AND2XL U_g249 (.A(G392GAT_23_gat), .B(G1GAT_0_gat), .Y(G564GAT_280_gat) );
AND2XL U_g250 (.A(G375GAT_22_gat), .B(G1GAT_0_gat), .Y(G561GAT_281_gat) );
AND2XL U_g251 (.A(G358GAT_21_gat), .B(G1GAT_0_gat), .Y(G558GAT_282_gat) );
AND2XL U_g252 (.A(G341GAT_20_gat), .B(G1GAT_0_gat), .Y(G555GAT_283_gat) );
AND2XL U_g253 (.A(G324GAT_19_gat), .B(G1GAT_0_gat), .Y(G552GAT_284_gat) );
AND2XL U_g254 (.A(G307GAT_18_gat), .B(G1GAT_0_gat), .Y(G549GAT_285_gat) );
AND2XL U_g255 (.A(G290GAT_17_gat), .B(G1GAT_0_gat), .Y(G546GAT_286_gat) );
AND2XL U_g256 (.A(G273GAT_16_gat), .B(G1GAT_0_gat), .Y(G545GAT_287_gat) );
BUFX20 U_g257 (.A(G1263GAT_47_gat), .Y(G1367GAT_288_gat) );
BUFX20 U_g258 (.A(G1215GAT_63_gat), .Y(G1363GAT_289_gat) );
BUFX20 U_g259 (.A(G1167GAT_79_gat), .Y(G1359GAT_290_gat) );
BUFX20 U_g260 (.A(G1119GAT_95_gat), .Y(G1355GAT_291_gat) );
BUFX20 U_g261 (.A(G1071GAT_111_gat), .Y(G1351GAT_292_gat) );
BUFX20 U_g262 (.A(G1023GAT_127_gat), .Y(G1347GAT_293_gat) );
BUFX20 U_g263 (.A(G975GAT_143_gat), .Y(G1343GAT_294_gat) );
BUFX20 U_g264 (.A(G927GAT_159_gat), .Y(G1339GAT_295_gat) );
BUFX20 U_g265 (.A(G879GAT_175_gat), .Y(G1335GAT_296_gat) );
BUFX20 U_g266 (.A(G831GAT_191_gat), .Y(G1331GAT_297_gat) );
BUFX20 U_g267 (.A(G783GAT_207_gat), .Y(G1327GAT_298_gat) );
BUFX20 U_g268 (.A(G735GAT_223_gat), .Y(G1323GAT_299_gat) );
BUFX20 U_g269 (.A(G687GAT_239_gat), .Y(G1319GAT_300_gat) );
BUFX20 U_g270 (.A(G639GAT_255_gat), .Y(G1315GAT_301_gat) );
BUFX20 U_g271 (.A(G591GAT_271_gat), .Y(G1311GAT_302_gat) );
BUFX20 U_g272 (.A(G1367GAT_288_gat), .Y(G1400GAT_303_gat) );
AND2XL U_g273 (.A(G1367GAT_288_ngat), .B(G1263GAT_47_ngat), .Y(G1399GAT_304_gat) );
BUFX20 U_g274 (.A(G1363GAT_289_gat), .Y(G1398GAT_305_gat) );
AND2XL U_g275 (.A(G1363GAT_289_ngat), .B(G1215GAT_63_ngat), .Y(G1397GAT_306_gat) );
BUFX20 U_g276 (.A(G1359GAT_290_gat), .Y(G1396GAT_307_gat) );
AND2XL U_g277 (.A(G1359GAT_290_ngat), .B(G1167GAT_79_ngat), .Y(G1395GAT_308_gat) );
BUFX20 U_g278 (.A(G1355GAT_291_gat), .Y(G1394GAT_309_gat) );
AND2XL U_g279 (.A(G1355GAT_291_ngat), .B(G1119GAT_95_ngat), .Y(G1393GAT_310_gat) );
BUFX20 U_g280 (.A(G1351GAT_292_gat), .Y(G1392GAT_311_gat) );
AND2XL U_g281 (.A(G1351GAT_292_ngat), .B(G1071GAT_111_ngat), .Y(G1391GAT_312_gat) );
BUFX20 U_g282 (.A(G1347GAT_293_gat), .Y(G1390GAT_313_gat) );
AND2XL U_g283 (.A(G1347GAT_293_ngat), .B(G1023GAT_127_ngat), .Y(G1389GAT_314_gat) );
BUFX20 U_g284 (.A(G1343GAT_294_gat), .Y(G1388GAT_315_gat) );
AND2XL U_g285 (.A(G1343GAT_294_ngat), .B(G975GAT_143_ngat), .Y(G1387GAT_316_gat) );
BUFX20 U_g286 (.A(G1339GAT_295_gat), .Y(G1386GAT_317_gat) );
AND2XL U_g287 (.A(G1339GAT_295_ngat), .B(G927GAT_159_ngat), .Y(G1385GAT_318_gat) );
BUFX20 U_g288 (.A(G1335GAT_296_gat), .Y(G1384GAT_319_gat) );
AND2XL U_g289 (.A(G1335GAT_296_ngat), .B(G879GAT_175_ngat), .Y(G1383GAT_320_gat) );
BUFX20 U_g290 (.A(G1331GAT_297_gat), .Y(G1382GAT_321_gat) );
AND2XL U_g291 (.A(G1331GAT_297_ngat), .B(G831GAT_191_ngat), .Y(G1381GAT_322_gat) );
BUFX20 U_g292 (.A(G1327GAT_298_gat), .Y(G1380GAT_323_gat) );
AND2XL U_g293 (.A(G1327GAT_298_ngat), .B(G783GAT_207_ngat), .Y(G1379GAT_324_gat) );
BUFX20 U_g294 (.A(G1323GAT_299_gat), .Y(G1378GAT_325_gat) );
AND2XL U_g295 (.A(G1323GAT_299_ngat), .B(G735GAT_223_ngat), .Y(G1377GAT_326_gat) );
BUFX20 U_g296 (.A(G1319GAT_300_gat), .Y(G1376GAT_327_gat) );
AND2XL U_g297 (.A(G1319GAT_300_ngat), .B(G687GAT_239_ngat), .Y(G1375GAT_328_gat) );
BUFX20 U_g298 (.A(G1315GAT_301_gat), .Y(G1374GAT_329_gat) );
AND2XL U_g299 (.A(G1315GAT_301_ngat), .B(G639GAT_255_ngat), .Y(G1373GAT_330_gat) );
BUFX20 U_g300 (.A(G1311GAT_302_gat), .Y(G1372GAT_331_gat) );
AND2XL U_g301 (.A(G1311GAT_302_ngat), .B(G591GAT_271_ngat), .Y(G1371GAT_332_gat) );
AND2XL U_g302 (.A(G1400GAT_303_ngat), .B(G1399GAT_304_ngat), .Y(G1443GAT_333_gat) );
AND2XL U_g303 (.A(G1398GAT_305_ngat), .B(G1397GAT_306_ngat), .Y(G1440GAT_334_gat) );
AND2XL U_g304 (.A(G1396GAT_307_ngat), .B(G1395GAT_308_ngat), .Y(G1437GAT_335_gat) );
AND2XL U_g305 (.A(G1394GAT_309_ngat), .B(G1393GAT_310_ngat), .Y(G1434GAT_336_gat) );
AND2XL U_g306 (.A(G1392GAT_311_ngat), .B(G1391GAT_312_ngat), .Y(G1431GAT_337_gat) );
AND2XL U_g307 (.A(G1390GAT_313_ngat), .B(G1389GAT_314_ngat), .Y(G1428GAT_338_gat) );
AND2XL U_g308 (.A(G1388GAT_315_ngat), .B(G1387GAT_316_ngat), .Y(G1425GAT_339_gat) );
AND2XL U_g309 (.A(G1386GAT_317_ngat), .B(G1385GAT_318_ngat), .Y(G1422GAT_340_gat) );
AND2XL U_g310 (.A(G1384GAT_319_ngat), .B(G1383GAT_320_ngat), .Y(G1419GAT_341_gat) );
AND2XL U_g311 (.A(G1382GAT_321_ngat), .B(G1381GAT_322_ngat), .Y(G1416GAT_342_gat) );
AND2XL U_g312 (.A(G1380GAT_323_ngat), .B(G1379GAT_324_ngat), .Y(G1413GAT_343_gat) );
AND2XL U_g313 (.A(G1378GAT_325_ngat), .B(G1377GAT_326_ngat), .Y(G1410GAT_344_gat) );
AND2XL U_g314 (.A(G1376GAT_327_ngat), .B(G1375GAT_328_ngat), .Y(G1407GAT_345_gat) );
AND2XL U_g315 (.A(G1374GAT_329_ngat), .B(G1373GAT_330_ngat), .Y(G1404GAT_346_gat) );
AND2XL U_g316 (.A(G1372GAT_331_ngat), .B(G1371GAT_332_ngat), .Y(G1401GAT_347_gat) );
AND2XL U_g317 (.A(G1218GAT_62_ngat), .B(G1443GAT_333_ngat), .Y(G1502GAT_348_gat) );
AND2XL U_g318 (.A(G1170GAT_78_ngat), .B(G1440GAT_334_ngat), .Y(G1498GAT_349_gat) );
AND2XL U_g319 (.A(G1122GAT_94_ngat), .B(G1437GAT_335_ngat), .Y(G1494GAT_350_gat) );
AND2XL U_g320 (.A(G1074GAT_110_ngat), .B(G1434GAT_336_ngat), .Y(G1490GAT_351_gat) );
AND2XL U_g321 (.A(G1026GAT_126_ngat), .B(G1431GAT_337_ngat), .Y(G1486GAT_352_gat) );
AND2XL U_g322 (.A(G978GAT_142_ngat), .B(G1428GAT_338_ngat), .Y(G1482GAT_353_gat) );
AND2XL U_g323 (.A(G930GAT_158_ngat), .B(G1425GAT_339_ngat), .Y(G1478GAT_354_gat) );
AND2XL U_g324 (.A(G882GAT_174_ngat), .B(G1422GAT_340_ngat), .Y(G1474GAT_355_gat) );
AND2XL U_g325 (.A(G834GAT_190_ngat), .B(G1419GAT_341_ngat), .Y(G1470GAT_356_gat) );
AND2XL U_g326 (.A(G786GAT_206_ngat), .B(G1416GAT_342_ngat), .Y(G1466GAT_357_gat) );
AND2XL U_g327 (.A(G738GAT_222_ngat), .B(G1413GAT_343_ngat), .Y(G1462GAT_358_gat) );
AND2XL U_g328 (.A(G690GAT_238_ngat), .B(G1410GAT_344_ngat), .Y(G1458GAT_359_gat) );
AND2XL U_g329 (.A(G642GAT_254_ngat), .B(G1407GAT_345_ngat), .Y(G1454GAT_360_gat) );
AND2XL U_g330 (.A(G594GAT_270_ngat), .B(G1404GAT_346_ngat), .Y(G1450GAT_361_gat) );
AND2XL U_g331 (.A(G546GAT_286_ngat), .B(G1401GAT_347_ngat), .Y(G1446GAT_362_gat) );
AND2XL U_g332 (.A(G1502GAT_348_ngat), .B(G1367GAT_288_ngat), .Y(G1578GAT_363_gat) );
AND2XL U_g333 (.A(G1502GAT_348_ngat), .B(G1443GAT_333_ngat), .Y(G1576GAT_364_gat) );
AND2XL U_g334 (.A(G1218GAT_62_ngat), .B(G1502GAT_348_ngat), .Y(G1577GAT_365_gat) );
AND2XL U_g335 (.A(G1498GAT_349_ngat), .B(G1363GAT_289_ngat), .Y(G1573GAT_366_gat) );
AND2XL U_g336 (.A(G1498GAT_349_ngat), .B(G1440GAT_334_ngat), .Y(G1571GAT_367_gat) );
AND2XL U_g337 (.A(G1170GAT_78_ngat), .B(G1498GAT_349_ngat), .Y(G1572GAT_368_gat) );
AND2XL U_g338 (.A(G1494GAT_350_ngat), .B(G1359GAT_290_ngat), .Y(G1568GAT_369_gat) );
AND2XL U_g339 (.A(G1494GAT_350_ngat), .B(G1437GAT_335_ngat), .Y(G1566GAT_370_gat) );
AND2XL U_g340 (.A(G1122GAT_94_ngat), .B(G1494GAT_350_ngat), .Y(G1567GAT_371_gat) );
AND2XL U_g341 (.A(G1490GAT_351_ngat), .B(G1355GAT_291_ngat), .Y(G1563GAT_372_gat) );
AND2XL U_g342 (.A(G1490GAT_351_ngat), .B(G1434GAT_336_ngat), .Y(G1561GAT_373_gat) );
AND2XL U_g343 (.A(G1074GAT_110_ngat), .B(G1490GAT_351_ngat), .Y(G1562GAT_374_gat) );
AND2XL U_g344 (.A(G1486GAT_352_ngat), .B(G1351GAT_292_ngat), .Y(G1558GAT_375_gat) );
AND2XL U_g345 (.A(G1486GAT_352_ngat), .B(G1431GAT_337_ngat), .Y(G1556GAT_376_gat) );
AND2XL U_g346 (.A(G1026GAT_126_ngat), .B(G1486GAT_352_ngat), .Y(G1557GAT_377_gat) );
AND2XL U_g347 (.A(G1482GAT_353_ngat), .B(G1347GAT_293_ngat), .Y(G1553GAT_378_gat) );
AND2XL U_g348 (.A(G1482GAT_353_ngat), .B(G1428GAT_338_ngat), .Y(G1551GAT_379_gat) );
AND2XL U_g349 (.A(G978GAT_142_ngat), .B(G1482GAT_353_ngat), .Y(G1552GAT_380_gat) );
AND2XL U_g350 (.A(G1478GAT_354_ngat), .B(G1343GAT_294_ngat), .Y(G1548GAT_381_gat) );
AND2XL U_g351 (.A(G1478GAT_354_ngat), .B(G1425GAT_339_ngat), .Y(G1546GAT_382_gat) );
AND2XL U_g352 (.A(G930GAT_158_ngat), .B(G1478GAT_354_ngat), .Y(G1547GAT_383_gat) );
AND2XL U_g353 (.A(G1474GAT_355_ngat), .B(G1339GAT_295_ngat), .Y(G1543GAT_384_gat) );
AND2XL U_g354 (.A(G1474GAT_355_ngat), .B(G1422GAT_340_ngat), .Y(G1541GAT_385_gat) );
AND2XL U_g355 (.A(G882GAT_174_ngat), .B(G1474GAT_355_ngat), .Y(G1542GAT_386_gat) );
AND2XL U_g356 (.A(G1470GAT_356_ngat), .B(G1335GAT_296_ngat), .Y(G1538GAT_387_gat) );
AND2XL U_g357 (.A(G1470GAT_356_ngat), .B(G1419GAT_341_ngat), .Y(G1536GAT_388_gat) );
AND2XL U_g358 (.A(G834GAT_190_ngat), .B(G1470GAT_356_ngat), .Y(G1537GAT_389_gat) );
AND2XL U_g359 (.A(G1466GAT_357_ngat), .B(G1331GAT_297_ngat), .Y(G1533GAT_390_gat) );
AND2XL U_g360 (.A(G1466GAT_357_ngat), .B(G1416GAT_342_ngat), .Y(G1531GAT_391_gat) );
AND2XL U_g361 (.A(G786GAT_206_ngat), .B(G1466GAT_357_ngat), .Y(G1532GAT_392_gat) );
AND2XL U_g362 (.A(G1462GAT_358_ngat), .B(G1327GAT_298_ngat), .Y(G1528GAT_393_gat) );
AND2XL U_g363 (.A(G1462GAT_358_ngat), .B(G1413GAT_343_ngat), .Y(G1526GAT_394_gat) );
AND2XL U_g364 (.A(G738GAT_222_ngat), .B(G1462GAT_358_ngat), .Y(G1527GAT_395_gat) );
AND2XL U_g365 (.A(G1458GAT_359_ngat), .B(G1323GAT_299_ngat), .Y(G1523GAT_396_gat) );
AND2XL U_g366 (.A(G1458GAT_359_ngat), .B(G1410GAT_344_ngat), .Y(G1521GAT_397_gat) );
AND2XL U_g367 (.A(G690GAT_238_ngat), .B(G1458GAT_359_ngat), .Y(G1522GAT_398_gat) );
AND2XL U_g368 (.A(G1454GAT_360_ngat), .B(G1319GAT_300_ngat), .Y(G1518GAT_399_gat) );
AND2XL U_g369 (.A(G1454GAT_360_ngat), .B(G1407GAT_345_ngat), .Y(G1516GAT_400_gat) );
AND2XL U_g370 (.A(G642GAT_254_ngat), .B(G1454GAT_360_ngat), .Y(G1517GAT_401_gat) );
AND2XL U_g371 (.A(G1450GAT_361_ngat), .B(G1315GAT_301_ngat), .Y(G1513GAT_402_gat) );
AND2XL U_g372 (.A(G1450GAT_361_ngat), .B(G1404GAT_346_ngat), .Y(G1511GAT_403_gat) );
AND2XL U_g373 (.A(G594GAT_270_ngat), .B(G1450GAT_361_ngat), .Y(G1512GAT_404_gat) );
AND2XL U_g374 (.A(G1446GAT_362_ngat), .B(G1311GAT_302_ngat), .Y(G1508GAT_405_gat) );
AND2XL U_g375 (.A(G1446GAT_362_ngat), .B(G1401GAT_347_ngat), .Y(G1506GAT_406_gat) );
AND2XL U_g376 (.A(G546GAT_286_ngat), .B(G1446GAT_362_ngat), .Y(G1507GAT_407_gat) );
AND2XL U_g377 (.A(G1578GAT_363_ngat), .B(G1266GAT_46_ngat), .Y(G1624GAT_408_gat) );
AND2XL U_g378 (.A(G1577GAT_365_ngat), .B(G1576GAT_364_ngat), .Y(G1621GAT_409_gat) );
AND2XL U_g379 (.A(G1572GAT_368_ngat), .B(G1571GAT_367_ngat), .Y(G1618GAT_410_gat) );
AND2XL U_g380 (.A(G1567GAT_371_ngat), .B(G1566GAT_370_ngat), .Y(G1615GAT_411_gat) );
AND2XL U_g381 (.A(G1562GAT_374_ngat), .B(G1561GAT_373_ngat), .Y(G1612GAT_412_gat) );
AND2XL U_g382 (.A(G1557GAT_377_ngat), .B(G1556GAT_376_ngat), .Y(G1609GAT_413_gat) );
AND2XL U_g383 (.A(G1552GAT_380_ngat), .B(G1551GAT_379_ngat), .Y(G1606GAT_414_gat) );
AND2XL U_g384 (.A(G1547GAT_383_ngat), .B(G1546GAT_382_ngat), .Y(G1603GAT_415_gat) );
AND2XL U_g385 (.A(G1542GAT_386_ngat), .B(G1541GAT_385_ngat), .Y(G1600GAT_416_gat) );
AND2XL U_g386 (.A(G1537GAT_389_ngat), .B(G1536GAT_388_ngat), .Y(G1597GAT_417_gat) );
AND2XL U_g387 (.A(G1532GAT_392_ngat), .B(G1531GAT_391_ngat), .Y(G1594GAT_418_gat) );
AND2XL U_g388 (.A(G1527GAT_395_ngat), .B(G1526GAT_394_ngat), .Y(G1591GAT_419_gat) );
AND2XL U_g389 (.A(G1522GAT_398_ngat), .B(G1521GAT_397_ngat), .Y(G1588GAT_420_gat) );
AND2XL U_g390 (.A(G1517GAT_401_ngat), .B(G1516GAT_400_ngat), .Y(G1585GAT_421_gat) );
AND2XL U_g391 (.A(G1512GAT_404_ngat), .B(G1511GAT_403_ngat), .Y(G1582GAT_422_gat) );
AND2XL U_g392 (.A(G1507GAT_407_ngat), .B(G1506GAT_406_ngat), .Y(G1581GAT_423_gat) );
AND2XL U_g393 (.A(G1624GAT_408_ngat), .B(G1266GAT_46_ngat), .Y(G1684GAT_424_gat) );
AND2XL U_g394 (.A(G1578GAT_363_ngat), .B(G1624GAT_408_ngat), .Y(G1685GAT_425_gat) );
AND2XL U_g395 (.A(G1573GAT_366_ngat), .B(G1621GAT_409_ngat), .Y(G1680GAT_426_gat) );
AND2XL U_g396 (.A(G1568GAT_369_ngat), .B(G1618GAT_410_ngat), .Y(G1676GAT_427_gat) );
AND2XL U_g397 (.A(G1563GAT_372_ngat), .B(G1615GAT_411_ngat), .Y(G1672GAT_428_gat) );
AND2XL U_g398 (.A(G1558GAT_375_ngat), .B(G1612GAT_412_ngat), .Y(G1668GAT_429_gat) );
AND2XL U_g399 (.A(G1553GAT_378_ngat), .B(G1609GAT_413_ngat), .Y(G1664GAT_430_gat) );
AND2XL U_g400 (.A(G1548GAT_381_ngat), .B(G1606GAT_414_ngat), .Y(G1660GAT_431_gat) );
AND2XL U_g401 (.A(G1543GAT_384_ngat), .B(G1603GAT_415_ngat), .Y(G1656GAT_432_gat) );
AND2XL U_g402 (.A(G1538GAT_387_ngat), .B(G1600GAT_416_ngat), .Y(G1652GAT_433_gat) );
AND2XL U_g403 (.A(G1533GAT_390_ngat), .B(G1597GAT_417_ngat), .Y(G1648GAT_434_gat) );
AND2XL U_g404 (.A(G1528GAT_393_ngat), .B(G1594GAT_418_ngat), .Y(G1644GAT_435_gat) );
AND2XL U_g405 (.A(G1523GAT_396_ngat), .B(G1591GAT_419_ngat), .Y(G1640GAT_436_gat) );
AND2XL U_g406 (.A(G1518GAT_399_ngat), .B(G1588GAT_420_ngat), .Y(G1636GAT_437_gat) );
AND2XL U_g407 (.A(G1513GAT_402_ngat), .B(G1585GAT_421_ngat), .Y(G1632GAT_438_gat) );
AND2XL U_g408 (.A(G1508GAT_405_ngat), .B(G1582GAT_422_ngat), .Y(G1628GAT_439_gat) );
AND2XL U_g409 (.A(G1685GAT_425_ngat), .B(G1684GAT_424_ngat), .Y(G1714GAT_440_gat) );
AND2XL U_g410 (.A(G1680GAT_426_ngat), .B(G1621GAT_409_ngat), .Y(G1712GAT_441_gat) );
AND2XL U_g411 (.A(G1573GAT_366_ngat), .B(G1680GAT_426_ngat), .Y(G1713GAT_442_gat) );
AND2XL U_g412 (.A(G1676GAT_427_ngat), .B(G1618GAT_410_ngat), .Y(G1710GAT_443_gat) );
AND2XL U_g413 (.A(G1568GAT_369_ngat), .B(G1676GAT_427_ngat), .Y(G1711GAT_444_gat) );
AND2XL U_g414 (.A(G1672GAT_428_ngat), .B(G1615GAT_411_ngat), .Y(G1708GAT_445_gat) );
AND2XL U_g415 (.A(G1563GAT_372_ngat), .B(G1672GAT_428_ngat), .Y(G1709GAT_446_gat) );
AND2XL U_g416 (.A(G1668GAT_429_ngat), .B(G1612GAT_412_ngat), .Y(G1706GAT_447_gat) );
AND2XL U_g417 (.A(G1558GAT_375_ngat), .B(G1668GAT_429_ngat), .Y(G1707GAT_448_gat) );
AND2XL U_g418 (.A(G1664GAT_430_ngat), .B(G1609GAT_413_ngat), .Y(G1704GAT_449_gat) );
AND2XL U_g419 (.A(G1553GAT_378_ngat), .B(G1664GAT_430_ngat), .Y(G1705GAT_450_gat) );
AND2XL U_g420 (.A(G1660GAT_431_ngat), .B(G1606GAT_414_ngat), .Y(G1702GAT_451_gat) );
AND2XL U_g421 (.A(G1548GAT_381_ngat), .B(G1660GAT_431_ngat), .Y(G1703GAT_452_gat) );
AND2XL U_g422 (.A(G1656GAT_432_ngat), .B(G1603GAT_415_ngat), .Y(G1700GAT_453_gat) );
AND2XL U_g423 (.A(G1543GAT_384_ngat), .B(G1656GAT_432_ngat), .Y(G1701GAT_454_gat) );
AND2XL U_g424 (.A(G1652GAT_433_ngat), .B(G1600GAT_416_ngat), .Y(G1698GAT_455_gat) );
AND2XL U_g425 (.A(G1538GAT_387_ngat), .B(G1652GAT_433_ngat), .Y(G1699GAT_456_gat) );
AND2XL U_g426 (.A(G1648GAT_434_ngat), .B(G1597GAT_417_ngat), .Y(G1696GAT_457_gat) );
AND2XL U_g427 (.A(G1533GAT_390_ngat), .B(G1648GAT_434_ngat), .Y(G1697GAT_458_gat) );
AND2XL U_g428 (.A(G1644GAT_435_ngat), .B(G1594GAT_418_ngat), .Y(G1694GAT_459_gat) );
AND2XL U_g429 (.A(G1528GAT_393_ngat), .B(G1644GAT_435_ngat), .Y(G1695GAT_460_gat) );
AND2XL U_g430 (.A(G1640GAT_436_ngat), .B(G1591GAT_419_ngat), .Y(G1692GAT_461_gat) );
AND2XL U_g431 (.A(G1523GAT_396_ngat), .B(G1640GAT_436_ngat), .Y(G1693GAT_462_gat) );
AND2XL U_g432 (.A(G1636GAT_437_ngat), .B(G1588GAT_420_ngat), .Y(G1690GAT_463_gat) );
AND2XL U_g433 (.A(G1518GAT_399_ngat), .B(G1636GAT_437_ngat), .Y(G1691GAT_464_gat) );
AND2XL U_g434 (.A(G1632GAT_438_ngat), .B(G1585GAT_421_ngat), .Y(G1688GAT_465_gat) );
AND2XL U_g435 (.A(G1513GAT_402_ngat), .B(G1632GAT_438_ngat), .Y(G1689GAT_466_gat) );
AND2XL U_g436 (.A(G1628GAT_439_ngat), .B(G1582GAT_422_ngat), .Y(G1686GAT_467_gat) );
AND2XL U_g437 (.A(G1508GAT_405_ngat), .B(G1628GAT_439_ngat), .Y(G1687GAT_468_gat) );
AND2XL U_g438 (.A(G1713GAT_442_ngat), .B(G1712GAT_441_ngat), .Y(G1756GAT_469_gat) );
AND2XL U_g439 (.A(G1221GAT_61_ngat), .B(G1714GAT_440_ngat), .Y(G1759GAT_470_gat) );
AND2XL U_g440 (.A(G1711GAT_444_ngat), .B(G1710GAT_443_ngat), .Y(G1753GAT_471_gat) );
AND2XL U_g441 (.A(G1709GAT_446_ngat), .B(G1708GAT_445_ngat), .Y(G1750GAT_472_gat) );
AND2XL U_g442 (.A(G1707GAT_448_ngat), .B(G1706GAT_447_ngat), .Y(G1747GAT_473_gat) );
AND2XL U_g443 (.A(G1705GAT_450_ngat), .B(G1704GAT_449_ngat), .Y(G1744GAT_474_gat) );
AND2XL U_g444 (.A(G1703GAT_452_ngat), .B(G1702GAT_451_ngat), .Y(G1741GAT_475_gat) );
AND2XL U_g445 (.A(G1701GAT_454_ngat), .B(G1700GAT_453_ngat), .Y(G1738GAT_476_gat) );
AND2XL U_g446 (.A(G1699GAT_456_ngat), .B(G1698GAT_455_ngat), .Y(G1735GAT_477_gat) );
AND2XL U_g447 (.A(G1697GAT_458_ngat), .B(G1696GAT_457_ngat), .Y(G1732GAT_478_gat) );
AND2XL U_g448 (.A(G1695GAT_460_ngat), .B(G1694GAT_459_ngat), .Y(G1729GAT_479_gat) );
AND2XL U_g449 (.A(G1693GAT_462_ngat), .B(G1692GAT_461_ngat), .Y(G1726GAT_480_gat) );
AND2XL U_g450 (.A(G1691GAT_464_ngat), .B(G1690GAT_463_ngat), .Y(G1723GAT_481_gat) );
AND2XL U_g451 (.A(G1689GAT_466_ngat), .B(G1688GAT_465_ngat), .Y(G1720GAT_482_gat) );
AND2XL U_g452 (.A(G1687GAT_468_ngat), .B(G1686GAT_467_ngat), .Y(G1717GAT_483_gat) );
AND2XL U_g453 (.A(G1759GAT_470_ngat), .B(G1624GAT_408_ngat), .Y(G1821GAT_484_gat) );
AND2XL U_g454 (.A(G1759GAT_470_ngat), .B(G1714GAT_440_ngat), .Y(G1819GAT_485_gat) );
AND2XL U_g455 (.A(G1221GAT_61_ngat), .B(G1759GAT_470_ngat), .Y(G1820GAT_486_gat) );
AND2XL U_g456 (.A(G1173GAT_77_ngat), .B(G1756GAT_469_ngat), .Y(G1815GAT_487_gat) );
AND2XL U_g457 (.A(G1125GAT_93_ngat), .B(G1753GAT_471_ngat), .Y(G1811GAT_488_gat) );
AND2XL U_g458 (.A(G1077GAT_109_ngat), .B(G1750GAT_472_ngat), .Y(G1807GAT_489_gat) );
AND2XL U_g459 (.A(G1029GAT_125_ngat), .B(G1747GAT_473_ngat), .Y(G1803GAT_490_gat) );
AND2XL U_g460 (.A(G981GAT_141_ngat), .B(G1744GAT_474_ngat), .Y(G1799GAT_491_gat) );
AND2XL U_g461 (.A(G933GAT_157_ngat), .B(G1741GAT_475_ngat), .Y(G1795GAT_492_gat) );
AND2XL U_g462 (.A(G885GAT_173_ngat), .B(G1738GAT_476_ngat), .Y(G1791GAT_493_gat) );
AND2XL U_g463 (.A(G837GAT_189_ngat), .B(G1735GAT_477_ngat), .Y(G1787GAT_494_gat) );
AND2XL U_g464 (.A(G789GAT_205_ngat), .B(G1732GAT_478_ngat), .Y(G1783GAT_495_gat) );
AND2XL U_g465 (.A(G741GAT_221_ngat), .B(G1729GAT_479_ngat), .Y(G1779GAT_496_gat) );
AND2XL U_g466 (.A(G693GAT_237_ngat), .B(G1726GAT_480_ngat), .Y(G1775GAT_497_gat) );
AND2XL U_g467 (.A(G645GAT_253_ngat), .B(G1723GAT_481_ngat), .Y(G1771GAT_498_gat) );
AND2XL U_g468 (.A(G597GAT_269_ngat), .B(G1720GAT_482_ngat), .Y(G1767GAT_499_gat) );
AND2XL U_g469 (.A(G549GAT_285_ngat), .B(G1717GAT_483_ngat), .Y(G1763GAT_500_gat) );
AND2XL U_g470 (.A(G1821GAT_484_ngat), .B(G1269GAT_45_ngat), .Y(G1897GAT_501_gat) );
AND2XL U_g471 (.A(G1820GAT_486_ngat), .B(G1819GAT_485_ngat), .Y(G1894GAT_502_gat) );
AND2XL U_g472 (.A(G1815GAT_487_ngat), .B(G1756GAT_469_ngat), .Y(G1889GAT_503_gat) );
AND2XL U_g473 (.A(G1815GAT_487_ngat), .B(G1680GAT_426_ngat), .Y(G1891GAT_504_gat) );
AND2XL U_g474 (.A(G1811GAT_488_ngat), .B(G1753GAT_471_ngat), .Y(G1884GAT_505_gat) );
AND2XL U_g475 (.A(G1173GAT_77_ngat), .B(G1815GAT_487_ngat), .Y(G1890GAT_506_gat) );
AND2XL U_g476 (.A(G1811GAT_488_ngat), .B(G1676GAT_427_ngat), .Y(G1886GAT_507_gat) );
AND2XL U_g477 (.A(G1807GAT_489_ngat), .B(G1750GAT_472_ngat), .Y(G1879GAT_508_gat) );
AND2XL U_g478 (.A(G1125GAT_93_ngat), .B(G1811GAT_488_ngat), .Y(G1885GAT_509_gat) );
AND2XL U_g479 (.A(G1807GAT_489_ngat), .B(G1672GAT_428_ngat), .Y(G1881GAT_510_gat) );
AND2XL U_g480 (.A(G1803GAT_490_ngat), .B(G1747GAT_473_ngat), .Y(G1874GAT_511_gat) );
AND2XL U_g481 (.A(G1077GAT_109_ngat), .B(G1807GAT_489_ngat), .Y(G1880GAT_512_gat) );
AND2XL U_g482 (.A(G1803GAT_490_ngat), .B(G1668GAT_429_ngat), .Y(G1876GAT_513_gat) );
AND2XL U_g483 (.A(G1799GAT_491_ngat), .B(G1744GAT_474_ngat), .Y(G1869GAT_514_gat) );
AND2XL U_g484 (.A(G1029GAT_125_ngat), .B(G1803GAT_490_ngat), .Y(G1875GAT_515_gat) );
AND2XL U_g485 (.A(G1799GAT_491_ngat), .B(G1664GAT_430_ngat), .Y(G1871GAT_516_gat) );
AND2XL U_g486 (.A(G1795GAT_492_ngat), .B(G1741GAT_475_ngat), .Y(G1864GAT_517_gat) );
AND2XL U_g487 (.A(G981GAT_141_ngat), .B(G1799GAT_491_ngat), .Y(G1870GAT_518_gat) );
AND2XL U_g488 (.A(G1795GAT_492_ngat), .B(G1660GAT_431_ngat), .Y(G1866GAT_519_gat) );
AND2XL U_g489 (.A(G1791GAT_493_ngat), .B(G1738GAT_476_ngat), .Y(G1859GAT_520_gat) );
AND2XL U_g490 (.A(G933GAT_157_ngat), .B(G1795GAT_492_ngat), .Y(G1865GAT_521_gat) );
AND2XL U_g491 (.A(G1791GAT_493_ngat), .B(G1656GAT_432_ngat), .Y(G1861GAT_522_gat) );
AND2XL U_g492 (.A(G1787GAT_494_ngat), .B(G1735GAT_477_ngat), .Y(G1854GAT_523_gat) );
AND2XL U_g493 (.A(G885GAT_173_ngat), .B(G1791GAT_493_ngat), .Y(G1860GAT_524_gat) );
AND2XL U_g494 (.A(G1787GAT_494_ngat), .B(G1652GAT_433_ngat), .Y(G1856GAT_525_gat) );
AND2XL U_g495 (.A(G1783GAT_495_ngat), .B(G1732GAT_478_ngat), .Y(G1849GAT_526_gat) );
AND2XL U_g496 (.A(G837GAT_189_ngat), .B(G1787GAT_494_ngat), .Y(G1855GAT_527_gat) );
AND2XL U_g497 (.A(G1783GAT_495_ngat), .B(G1648GAT_434_ngat), .Y(G1851GAT_528_gat) );
AND2XL U_g498 (.A(G1779GAT_496_ngat), .B(G1729GAT_479_ngat), .Y(G1844GAT_529_gat) );
AND2XL U_g499 (.A(G789GAT_205_ngat), .B(G1783GAT_495_ngat), .Y(G1850GAT_530_gat) );
AND2XL U_g500 (.A(G1779GAT_496_ngat), .B(G1644GAT_435_ngat), .Y(G1846GAT_531_gat) );
AND2XL U_g501 (.A(G1775GAT_497_ngat), .B(G1726GAT_480_ngat), .Y(G1839GAT_532_gat) );
AND2XL U_g502 (.A(G741GAT_221_ngat), .B(G1779GAT_496_ngat), .Y(G1845GAT_533_gat) );
AND2XL U_g503 (.A(G1775GAT_497_ngat), .B(G1640GAT_436_ngat), .Y(G1841GAT_534_gat) );
AND2XL U_g504 (.A(G1771GAT_498_ngat), .B(G1723GAT_481_ngat), .Y(G1834GAT_535_gat) );
AND2XL U_g505 (.A(G693GAT_237_ngat), .B(G1775GAT_497_ngat), .Y(G1840GAT_536_gat) );
AND2XL U_g506 (.A(G1771GAT_498_ngat), .B(G1636GAT_437_ngat), .Y(G1836GAT_537_gat) );
AND2XL U_g507 (.A(G1767GAT_499_ngat), .B(G1720GAT_482_ngat), .Y(G1829GAT_538_gat) );
AND2XL U_g508 (.A(G645GAT_253_ngat), .B(G1771GAT_498_ngat), .Y(G1835GAT_539_gat) );
AND2XL U_g509 (.A(G1767GAT_499_ngat), .B(G1632GAT_438_ngat), .Y(G1831GAT_540_gat) );
AND2XL U_g510 (.A(G1763GAT_500_ngat), .B(G1717GAT_483_ngat), .Y(G1824GAT_541_gat) );
AND2XL U_g511 (.A(G597GAT_269_ngat), .B(G1767GAT_499_ngat), .Y(G1830GAT_542_gat) );
AND2XL U_g512 (.A(G1763GAT_500_ngat), .B(G1628GAT_439_ngat), .Y(G1826GAT_543_gat) );
AND2XL U_g513 (.A(G549GAT_285_ngat), .B(G1763GAT_500_ngat), .Y(G1825GAT_544_gat) );
AND2XL U_g514 (.A(G1897GAT_501_ngat), .B(G1269GAT_45_ngat), .Y(G1945GAT_545_gat) );
AND2XL U_g515 (.A(G1821GAT_484_ngat), .B(G1897GAT_501_ngat), .Y(G1946GAT_546_gat) );
AND2XL U_g516 (.A(G1891GAT_504_ngat), .B(G1894GAT_502_ngat), .Y(G1941GAT_547_gat) );
AND2XL U_g517 (.A(G1890GAT_506_ngat), .B(G1889GAT_503_ngat), .Y(G1938GAT_548_gat) );
AND2XL U_g518 (.A(G1885GAT_509_ngat), .B(G1884GAT_505_ngat), .Y(G1935GAT_549_gat) );
AND2XL U_g519 (.A(G1880GAT_512_ngat), .B(G1879GAT_508_ngat), .Y(G1932GAT_550_gat) );
AND2XL U_g520 (.A(G1875GAT_515_ngat), .B(G1874GAT_511_ngat), .Y(G1929GAT_551_gat) );
AND2XL U_g521 (.A(G1870GAT_518_ngat), .B(G1869GAT_514_ngat), .Y(G1926GAT_552_gat) );
AND2XL U_g522 (.A(G1865GAT_521_ngat), .B(G1864GAT_517_ngat), .Y(G1923GAT_553_gat) );
AND2XL U_g523 (.A(G1860GAT_524_ngat), .B(G1859GAT_520_ngat), .Y(G1920GAT_554_gat) );
AND2XL U_g524 (.A(G1855GAT_527_ngat), .B(G1854GAT_523_ngat), .Y(G1917GAT_555_gat) );
AND2XL U_g525 (.A(G1850GAT_530_ngat), .B(G1849GAT_526_ngat), .Y(G1914GAT_556_gat) );
AND2XL U_g526 (.A(G1845GAT_533_ngat), .B(G1844GAT_529_ngat), .Y(G1911GAT_557_gat) );
AND2XL U_g527 (.A(G1840GAT_536_ngat), .B(G1839GAT_532_ngat), .Y(G1908GAT_558_gat) );
AND2XL U_g528 (.A(G1835GAT_539_ngat), .B(G1834GAT_535_ngat), .Y(G1905GAT_559_gat) );
AND2XL U_g529 (.A(G1830GAT_542_ngat), .B(G1829GAT_538_ngat), .Y(G1902GAT_560_gat) );
AND2XL U_g530 (.A(G1825GAT_544_ngat), .B(G1824GAT_541_ngat), .Y(G1901GAT_561_gat) );
AND2XL U_g531 (.A(G1946GAT_546_ngat), .B(G1945GAT_545_ngat), .Y(G2001GAT_562_gat) );
AND2XL U_g532 (.A(G1941GAT_547_ngat), .B(G1894GAT_502_ngat), .Y(G1999GAT_563_gat) );
AND2XL U_g533 (.A(G1891GAT_504_ngat), .B(G1941GAT_547_ngat), .Y(G2000GAT_564_gat) );
AND2XL U_g534 (.A(G1886GAT_507_ngat), .B(G1938GAT_548_ngat), .Y(G1995GAT_565_gat) );
AND2XL U_g535 (.A(G1881GAT_510_ngat), .B(G1935GAT_549_ngat), .Y(G1991GAT_566_gat) );
AND2XL U_g536 (.A(G1876GAT_513_ngat), .B(G1932GAT_550_ngat), .Y(G1987GAT_567_gat) );
AND2XL U_g537 (.A(G1871GAT_516_ngat), .B(G1929GAT_551_ngat), .Y(G1983GAT_568_gat) );
AND2XL U_g538 (.A(G1866GAT_519_ngat), .B(G1926GAT_552_ngat), .Y(G1979GAT_569_gat) );
AND2XL U_g539 (.A(G1861GAT_522_ngat), .B(G1923GAT_553_ngat), .Y(G1975GAT_570_gat) );
AND2XL U_g540 (.A(G1856GAT_525_ngat), .B(G1920GAT_554_ngat), .Y(G1971GAT_571_gat) );
AND2XL U_g541 (.A(G1851GAT_528_ngat), .B(G1917GAT_555_ngat), .Y(G1967GAT_572_gat) );
AND2XL U_g542 (.A(G1846GAT_531_ngat), .B(G1914GAT_556_ngat), .Y(G1963GAT_573_gat) );
AND2XL U_g543 (.A(G1841GAT_534_ngat), .B(G1911GAT_557_ngat), .Y(G1959GAT_574_gat) );
AND2XL U_g544 (.A(G1836GAT_537_ngat), .B(G1908GAT_558_ngat), .Y(G1955GAT_575_gat) );
AND2XL U_g545 (.A(G1831GAT_540_ngat), .B(G1905GAT_559_ngat), .Y(G1951GAT_576_gat) );
AND2XL U_g546 (.A(G1826GAT_543_ngat), .B(G1902GAT_560_ngat), .Y(G1947GAT_577_gat) );
AND2XL U_g547 (.A(G2000GAT_564_ngat), .B(G1999GAT_563_ngat), .Y(G2030GAT_578_gat) );
AND2XL U_g548 (.A(G1995GAT_565_ngat), .B(G1938GAT_548_ngat), .Y(G2028GAT_579_gat) );
AND2XL U_g549 (.A(G1224GAT_60_ngat), .B(G2001GAT_562_ngat), .Y(G2033GAT_580_gat) );
AND2XL U_g550 (.A(G1991GAT_566_ngat), .B(G1935GAT_549_ngat), .Y(G2026GAT_581_gat) );
AND2XL U_g551 (.A(G1886GAT_507_ngat), .B(G1995GAT_565_ngat), .Y(G2029GAT_582_gat) );
AND2XL U_g552 (.A(G1987GAT_567_ngat), .B(G1932GAT_550_ngat), .Y(G2024GAT_583_gat) );
AND2XL U_g553 (.A(G1881GAT_510_ngat), .B(G1991GAT_566_ngat), .Y(G2027GAT_584_gat) );
AND2XL U_g554 (.A(G1983GAT_568_ngat), .B(G1929GAT_551_ngat), .Y(G2022GAT_585_gat) );
AND2XL U_g555 (.A(G1876GAT_513_ngat), .B(G1987GAT_567_ngat), .Y(G2025GAT_586_gat) );
AND2XL U_g556 (.A(G1979GAT_569_ngat), .B(G1926GAT_552_ngat), .Y(G2020GAT_587_gat) );
AND2XL U_g557 (.A(G1871GAT_516_ngat), .B(G1983GAT_568_ngat), .Y(G2023GAT_588_gat) );
AND2XL U_g558 (.A(G1975GAT_570_ngat), .B(G1923GAT_553_ngat), .Y(G2018GAT_589_gat) );
AND2XL U_g559 (.A(G1866GAT_519_ngat), .B(G1979GAT_569_ngat), .Y(G2021GAT_590_gat) );
AND2XL U_g560 (.A(G1971GAT_571_ngat), .B(G1920GAT_554_ngat), .Y(G2016GAT_591_gat) );
AND2XL U_g561 (.A(G1861GAT_522_ngat), .B(G1975GAT_570_ngat), .Y(G2019GAT_592_gat) );
AND2XL U_g562 (.A(G1967GAT_572_ngat), .B(G1917GAT_555_ngat), .Y(G2014GAT_593_gat) );
AND2XL U_g563 (.A(G1856GAT_525_ngat), .B(G1971GAT_571_ngat), .Y(G2017GAT_594_gat) );
AND2XL U_g564 (.A(G1963GAT_573_ngat), .B(G1914GAT_556_ngat), .Y(G2012GAT_595_gat) );
AND2XL U_g565 (.A(G1851GAT_528_ngat), .B(G1967GAT_572_ngat), .Y(G2015GAT_596_gat) );
AND2XL U_g566 (.A(G1959GAT_574_ngat), .B(G1911GAT_557_ngat), .Y(G2010GAT_597_gat) );
AND2XL U_g567 (.A(G1846GAT_531_ngat), .B(G1963GAT_573_ngat), .Y(G2013GAT_598_gat) );
AND2XL U_g568 (.A(G1955GAT_575_ngat), .B(G1908GAT_558_ngat), .Y(G2008GAT_599_gat) );
AND2XL U_g569 (.A(G1841GAT_534_ngat), .B(G1959GAT_574_ngat), .Y(G2011GAT_600_gat) );
AND2XL U_g570 (.A(G1951GAT_576_ngat), .B(G1905GAT_559_ngat), .Y(G2006GAT_601_gat) );
AND2XL U_g571 (.A(G1836GAT_537_ngat), .B(G1955GAT_575_ngat), .Y(G2009GAT_602_gat) );
AND2XL U_g572 (.A(G1947GAT_577_ngat), .B(G1902GAT_560_ngat), .Y(G2004GAT_603_gat) );
AND2XL U_g573 (.A(G1831GAT_540_ngat), .B(G1951GAT_576_ngat), .Y(G2007GAT_604_gat) );
AND2XL U_g574 (.A(G1826GAT_543_ngat), .B(G1947GAT_577_ngat), .Y(G2005GAT_605_gat) );
AND2XL U_g575 (.A(G2033GAT_580_ngat), .B(G1897GAT_501_ngat), .Y(G2082GAT_606_gat) );
AND2XL U_g576 (.A(G2033GAT_580_ngat), .B(G2001GAT_562_ngat), .Y(G2080GAT_607_gat) );
AND2XL U_g577 (.A(G2029GAT_582_ngat), .B(G2028GAT_579_ngat), .Y(G2073GAT_608_gat) );
AND2XL U_g578 (.A(G1224GAT_60_ngat), .B(G2033GAT_580_ngat), .Y(G2081GAT_609_gat) );
AND2XL U_g579 (.A(G2027GAT_584_ngat), .B(G2026GAT_581_ngat), .Y(G2070GAT_610_gat) );
AND2XL U_g580 (.A(G1176GAT_76_ngat), .B(G2030GAT_578_ngat), .Y(G2076GAT_611_gat) );
AND2XL U_g581 (.A(G2025GAT_586_ngat), .B(G2024GAT_583_ngat), .Y(G2067GAT_612_gat) );
AND2XL U_g582 (.A(G2023GAT_588_ngat), .B(G2022GAT_585_ngat), .Y(G2064GAT_613_gat) );
AND2XL U_g583 (.A(G2021GAT_590_ngat), .B(G2020GAT_587_ngat), .Y(G2061GAT_614_gat) );
AND2XL U_g584 (.A(G2019GAT_592_ngat), .B(G2018GAT_589_ngat), .Y(G2058GAT_615_gat) );
AND2XL U_g585 (.A(G2017GAT_594_ngat), .B(G2016GAT_591_ngat), .Y(G2055GAT_616_gat) );
AND2XL U_g586 (.A(G2015GAT_596_ngat), .B(G2014GAT_593_ngat), .Y(G2052GAT_617_gat) );
AND2XL U_g587 (.A(G2013GAT_598_ngat), .B(G2012GAT_595_ngat), .Y(G2049GAT_618_gat) );
AND2XL U_g588 (.A(G2011GAT_600_ngat), .B(G2010GAT_597_ngat), .Y(G2046GAT_619_gat) );
AND2XL U_g589 (.A(G2009GAT_602_ngat), .B(G2008GAT_599_ngat), .Y(G2043GAT_620_gat) );
AND2XL U_g590 (.A(G2007GAT_604_ngat), .B(G2006GAT_601_ngat), .Y(G2040GAT_621_gat) );
AND2XL U_g591 (.A(G2005GAT_605_ngat), .B(G2004GAT_603_ngat), .Y(G2037GAT_622_gat) );
AND2XL U_g592 (.A(G2082GAT_606_ngat), .B(G1272GAT_44_ngat), .Y(G2145GAT_623_gat) );
AND2XL U_g593 (.A(G2081GAT_609_ngat), .B(G2080GAT_607_ngat), .Y(G2142GAT_624_gat) );
AND2XL U_g594 (.A(G2076GAT_611_ngat), .B(G1941GAT_547_ngat), .Y(G2139GAT_625_gat) );
AND2XL U_g595 (.A(G2076GAT_611_ngat), .B(G2030GAT_578_ngat), .Y(G2137GAT_626_gat) );
AND2XL U_g596 (.A(G1176GAT_76_ngat), .B(G2076GAT_611_ngat), .Y(G2138GAT_627_gat) );
AND2XL U_g597 (.A(G1128GAT_92_ngat), .B(G2073GAT_608_ngat), .Y(G2133GAT_628_gat) );
AND2XL U_g598 (.A(G1080GAT_108_ngat), .B(G2070GAT_610_ngat), .Y(G2129GAT_629_gat) );
AND2XL U_g599 (.A(G1032GAT_124_ngat), .B(G2067GAT_612_ngat), .Y(G2125GAT_630_gat) );
AND2XL U_g600 (.A(G984GAT_140_ngat), .B(G2064GAT_613_ngat), .Y(G2121GAT_631_gat) );
AND2XL U_g601 (.A(G936GAT_156_ngat), .B(G2061GAT_614_ngat), .Y(G2117GAT_632_gat) );
AND2XL U_g602 (.A(G888GAT_172_ngat), .B(G2058GAT_615_ngat), .Y(G2113GAT_633_gat) );
AND2XL U_g603 (.A(G840GAT_188_ngat), .B(G2055GAT_616_ngat), .Y(G2109GAT_634_gat) );
AND2XL U_g604 (.A(G792GAT_204_ngat), .B(G2052GAT_617_ngat), .Y(G2105GAT_635_gat) );
AND2XL U_g605 (.A(G744GAT_220_ngat), .B(G2049GAT_618_ngat), .Y(G2101GAT_636_gat) );
AND2XL U_g606 (.A(G696GAT_236_ngat), .B(G2046GAT_619_ngat), .Y(G2097GAT_637_gat) );
AND2XL U_g607 (.A(G648GAT_252_ngat), .B(G2043GAT_620_ngat), .Y(G2093GAT_638_gat) );
AND2XL U_g608 (.A(G600GAT_268_ngat), .B(G2040GAT_621_ngat), .Y(G2089GAT_639_gat) );
AND2XL U_g609 (.A(G552GAT_284_ngat), .B(G2037GAT_622_ngat), .Y(G2085GAT_640_gat) );
AND2XL U_g610 (.A(G2145GAT_623_ngat), .B(G1272GAT_44_ngat), .Y(G2221GAT_641_gat) );
AND2XL U_g611 (.A(G2082GAT_606_ngat), .B(G2145GAT_623_ngat), .Y(G2222GAT_642_gat) );
AND2XL U_g612 (.A(G2139GAT_625_ngat), .B(G2142GAT_624_ngat), .Y(G2217GAT_643_gat) );
AND2XL U_g613 (.A(G2138GAT_627_ngat), .B(G2137GAT_626_ngat), .Y(G2214GAT_644_gat) );
AND2XL U_g614 (.A(G2133GAT_628_ngat), .B(G2073GAT_608_ngat), .Y(G2209GAT_645_gat) );
AND2XL U_g615 (.A(G2129GAT_629_ngat), .B(G2070GAT_610_ngat), .Y(G2204GAT_646_gat) );
AND2XL U_g616 (.A(G2133GAT_628_ngat), .B(G1995GAT_565_ngat), .Y(G2211GAT_647_gat) );
AND2XL U_g617 (.A(G2125GAT_630_ngat), .B(G2067GAT_612_ngat), .Y(G2199GAT_648_gat) );
AND2XL U_g618 (.A(G1128GAT_92_ngat), .B(G2133GAT_628_ngat), .Y(G2210GAT_649_gat) );
AND2XL U_g619 (.A(G2129GAT_629_ngat), .B(G1991GAT_566_ngat), .Y(G2206GAT_650_gat) );
AND2XL U_g620 (.A(G2121GAT_631_ngat), .B(G2064GAT_613_ngat), .Y(G2194GAT_651_gat) );
AND2XL U_g621 (.A(G1080GAT_108_ngat), .B(G2129GAT_629_ngat), .Y(G2205GAT_652_gat) );
AND2XL U_g622 (.A(G2125GAT_630_ngat), .B(G1987GAT_567_ngat), .Y(G2201GAT_653_gat) );
AND2XL U_g623 (.A(G2117GAT_632_ngat), .B(G2061GAT_614_ngat), .Y(G2189GAT_654_gat) );
AND2XL U_g624 (.A(G1032GAT_124_ngat), .B(G2125GAT_630_ngat), .Y(G2200GAT_655_gat) );
AND2XL U_g625 (.A(G2121GAT_631_ngat), .B(G1983GAT_568_ngat), .Y(G2196GAT_656_gat) );
AND2XL U_g626 (.A(G2113GAT_633_ngat), .B(G2058GAT_615_ngat), .Y(G2184GAT_657_gat) );
AND2XL U_g627 (.A(G984GAT_140_ngat), .B(G2121GAT_631_ngat), .Y(G2195GAT_658_gat) );
AND2XL U_g628 (.A(G2117GAT_632_ngat), .B(G1979GAT_569_ngat), .Y(G2191GAT_659_gat) );
AND2XL U_g629 (.A(G2109GAT_634_ngat), .B(G2055GAT_616_ngat), .Y(G2179GAT_660_gat) );
AND2XL U_g630 (.A(G936GAT_156_ngat), .B(G2117GAT_632_ngat), .Y(G2190GAT_661_gat) );
AND2XL U_g631 (.A(G2113GAT_633_ngat), .B(G1975GAT_570_ngat), .Y(G2186GAT_662_gat) );
AND2XL U_g632 (.A(G2105GAT_635_ngat), .B(G2052GAT_617_ngat), .Y(G2174GAT_663_gat) );
AND2XL U_g633 (.A(G888GAT_172_ngat), .B(G2113GAT_633_ngat), .Y(G2185GAT_664_gat) );
AND2XL U_g634 (.A(G2109GAT_634_ngat), .B(G1971GAT_571_ngat), .Y(G2181GAT_665_gat) );
AND2XL U_g635 (.A(G2101GAT_636_ngat), .B(G2049GAT_618_ngat), .Y(G2169GAT_666_gat) );
AND2XL U_g636 (.A(G840GAT_188_ngat), .B(G2109GAT_634_ngat), .Y(G2180GAT_667_gat) );
AND2XL U_g637 (.A(G2105GAT_635_ngat), .B(G1967GAT_572_ngat), .Y(G2176GAT_668_gat) );
AND2XL U_g638 (.A(G2097GAT_637_ngat), .B(G2046GAT_619_ngat), .Y(G2164GAT_669_gat) );
AND2XL U_g639 (.A(G792GAT_204_ngat), .B(G2105GAT_635_ngat), .Y(G2175GAT_670_gat) );
AND2XL U_g640 (.A(G2101GAT_636_ngat), .B(G1963GAT_573_ngat), .Y(G2171GAT_671_gat) );
AND2XL U_g641 (.A(G2093GAT_638_ngat), .B(G2043GAT_620_ngat), .Y(G2159GAT_672_gat) );
AND2XL U_g642 (.A(G744GAT_220_ngat), .B(G2101GAT_636_ngat), .Y(G2170GAT_673_gat) );
AND2XL U_g643 (.A(G2097GAT_637_ngat), .B(G1959GAT_574_ngat), .Y(G2166GAT_674_gat) );
AND2XL U_g644 (.A(G2089GAT_639_ngat), .B(G2040GAT_621_ngat), .Y(G2154GAT_675_gat) );
AND2XL U_g645 (.A(G696GAT_236_ngat), .B(G2097GAT_637_ngat), .Y(G2165GAT_676_gat) );
AND2XL U_g646 (.A(G2093GAT_638_ngat), .B(G1955GAT_575_ngat), .Y(G2161GAT_677_gat) );
AND2XL U_g647 (.A(G2085GAT_640_ngat), .B(G2037GAT_622_ngat), .Y(G2149GAT_678_gat) );
AND2XL U_g648 (.A(G648GAT_252_ngat), .B(G2093GAT_638_ngat), .Y(G2160GAT_679_gat) );
AND2XL U_g649 (.A(G2089GAT_639_ngat), .B(G1951GAT_576_ngat), .Y(G2156GAT_680_gat) );
AND2XL U_g650 (.A(G600GAT_268_ngat), .B(G2089GAT_639_ngat), .Y(G2155GAT_681_gat) );
AND2XL U_g651 (.A(G2085GAT_640_ngat), .B(G1947GAT_577_ngat), .Y(G2151GAT_682_gat) );
AND2XL U_g652 (.A(G552GAT_284_ngat), .B(G2085GAT_640_ngat), .Y(G2150GAT_683_gat) );
AND2XL U_g653 (.A(G2222GAT_642_ngat), .B(G2221GAT_641_ngat), .Y(G2266GAT_684_gat) );
AND2XL U_g654 (.A(G2217GAT_643_ngat), .B(G2142GAT_624_ngat), .Y(G2264GAT_685_gat) );
AND2XL U_g655 (.A(G2139GAT_625_ngat), .B(G2217GAT_643_ngat), .Y(G2265GAT_686_gat) );
AND2XL U_g656 (.A(G2211GAT_647_ngat), .B(G2214GAT_644_ngat), .Y(G2260GAT_687_gat) );
AND2XL U_g657 (.A(G2210GAT_649_ngat), .B(G2209GAT_645_ngat), .Y(G2257GAT_688_gat) );
AND2XL U_g658 (.A(G2205GAT_652_ngat), .B(G2204GAT_646_ngat), .Y(G2254GAT_689_gat) );
AND2XL U_g659 (.A(G2200GAT_655_ngat), .B(G2199GAT_648_ngat), .Y(G2251GAT_690_gat) );
AND2XL U_g660 (.A(G2195GAT_658_ngat), .B(G2194GAT_651_ngat), .Y(G2248GAT_691_gat) );
AND2XL U_g661 (.A(G2190GAT_661_ngat), .B(G2189GAT_654_ngat), .Y(G2245GAT_692_gat) );
AND2XL U_g662 (.A(G2185GAT_664_ngat), .B(G2184GAT_657_ngat), .Y(G2242GAT_693_gat) );
AND2XL U_g663 (.A(G2180GAT_667_ngat), .B(G2179GAT_660_ngat), .Y(G2239GAT_694_gat) );
AND2XL U_g664 (.A(G2175GAT_670_ngat), .B(G2174GAT_663_ngat), .Y(G2236GAT_695_gat) );
AND2XL U_g665 (.A(G2170GAT_673_ngat), .B(G2169GAT_666_ngat), .Y(G2233GAT_696_gat) );
AND2XL U_g666 (.A(G2165GAT_676_ngat), .B(G2164GAT_669_ngat), .Y(G2230GAT_697_gat) );
AND2XL U_g667 (.A(G2160GAT_679_ngat), .B(G2159GAT_672_ngat), .Y(G2227GAT_698_gat) );
AND2XL U_g668 (.A(G2155GAT_681_ngat), .B(G2154GAT_675_ngat), .Y(G2224GAT_699_gat) );
AND2XL U_g669 (.A(G2150GAT_683_ngat), .B(G2149GAT_678_ngat), .Y(G2223GAT_700_gat) );
AND2XL U_g670 (.A(G2265GAT_686_ngat), .B(G2264GAT_685_ngat), .Y(G2319GAT_701_gat) );
AND2XL U_g671 (.A(G2260GAT_687_ngat), .B(G2214GAT_644_ngat), .Y(G2317GAT_702_gat) );
AND2XL U_g672 (.A(G1227GAT_59_ngat), .B(G2266GAT_684_ngat), .Y(G2322GAT_703_gat) );
AND2XL U_g673 (.A(G2211GAT_647_ngat), .B(G2260GAT_687_ngat), .Y(G2318GAT_704_gat) );
AND2XL U_g674 (.A(G2206GAT_650_ngat), .B(G2257GAT_688_ngat), .Y(G2313GAT_705_gat) );
AND2XL U_g675 (.A(G2201GAT_653_ngat), .B(G2254GAT_689_ngat), .Y(G2309GAT_706_gat) );
AND2XL U_g676 (.A(G2196GAT_656_ngat), .B(G2251GAT_690_ngat), .Y(G2305GAT_707_gat) );
AND2XL U_g677 (.A(G2191GAT_659_ngat), .B(G2248GAT_691_ngat), .Y(G2301GAT_708_gat) );
AND2XL U_g678 (.A(G2186GAT_662_ngat), .B(G2245GAT_692_ngat), .Y(G2297GAT_709_gat) );
AND2XL U_g679 (.A(G2181GAT_665_ngat), .B(G2242GAT_693_ngat), .Y(G2293GAT_710_gat) );
AND2XL U_g680 (.A(G2176GAT_668_ngat), .B(G2239GAT_694_ngat), .Y(G2289GAT_711_gat) );
AND2XL U_g681 (.A(G2171GAT_671_ngat), .B(G2236GAT_695_ngat), .Y(G2285GAT_712_gat) );
AND2XL U_g682 (.A(G2166GAT_674_ngat), .B(G2233GAT_696_ngat), .Y(G2281GAT_713_gat) );
AND2XL U_g683 (.A(G2161GAT_677_ngat), .B(G2230GAT_697_ngat), .Y(G2277GAT_714_gat) );
AND2XL U_g684 (.A(G2156GAT_680_ngat), .B(G2227GAT_698_ngat), .Y(G2273GAT_715_gat) );
AND2XL U_g685 (.A(G2151GAT_682_ngat), .B(G2224GAT_699_ngat), .Y(G2269GAT_716_gat) );
AND2XL U_g686 (.A(G2322GAT_703_ngat), .B(G2145GAT_623_ngat), .Y(G2359GAT_717_gat) );
AND2XL U_g687 (.A(G2322GAT_703_ngat), .B(G2266GAT_684_ngat), .Y(G2357GAT_718_gat) );
AND2XL U_g688 (.A(G2318GAT_704_ngat), .B(G2317GAT_702_ngat), .Y(G2350GAT_719_gat) );
AND2XL U_g689 (.A(G2313GAT_705_ngat), .B(G2257GAT_688_ngat), .Y(G2348GAT_720_gat) );
AND2XL U_g690 (.A(G1227GAT_59_ngat), .B(G2322GAT_703_ngat), .Y(G2358GAT_721_gat) );
AND2XL U_g691 (.A(G2309GAT_706_ngat), .B(G2254GAT_689_ngat), .Y(G2346GAT_722_gat) );
AND2XL U_g692 (.A(G1179GAT_75_ngat), .B(G2319GAT_701_ngat), .Y(G2353GAT_723_gat) );
AND2XL U_g693 (.A(G2305GAT_707_ngat), .B(G2251GAT_690_ngat), .Y(G2344GAT_724_gat) );
AND2XL U_g694 (.A(G2206GAT_650_ngat), .B(G2313GAT_705_ngat), .Y(G2349GAT_725_gat) );
AND2XL U_g695 (.A(G2301GAT_708_ngat), .B(G2248GAT_691_ngat), .Y(G2342GAT_726_gat) );
AND2XL U_g696 (.A(G2201GAT_653_ngat), .B(G2309GAT_706_ngat), .Y(G2347GAT_727_gat) );
AND2XL U_g697 (.A(G2297GAT_709_ngat), .B(G2245GAT_692_ngat), .Y(G2340GAT_728_gat) );
AND2XL U_g698 (.A(G2196GAT_656_ngat), .B(G2305GAT_707_ngat), .Y(G2345GAT_729_gat) );
AND2XL U_g699 (.A(G2293GAT_710_ngat), .B(G2242GAT_693_ngat), .Y(G2338GAT_730_gat) );
AND2XL U_g700 (.A(G2191GAT_659_ngat), .B(G2301GAT_708_ngat), .Y(G2343GAT_731_gat) );
AND2XL U_g701 (.A(G2289GAT_711_ngat), .B(G2239GAT_694_ngat), .Y(G2336GAT_732_gat) );
AND2XL U_g702 (.A(G2186GAT_662_ngat), .B(G2297GAT_709_ngat), .Y(G2341GAT_733_gat) );
AND2XL U_g703 (.A(G2285GAT_712_ngat), .B(G2236GAT_695_ngat), .Y(G2334GAT_734_gat) );
AND2XL U_g704 (.A(G2181GAT_665_ngat), .B(G2293GAT_710_ngat), .Y(G2339GAT_735_gat) );
AND2XL U_g705 (.A(G2281GAT_713_ngat), .B(G2233GAT_696_ngat), .Y(G2332GAT_736_gat) );
AND2XL U_g706 (.A(G2176GAT_668_ngat), .B(G2289GAT_711_ngat), .Y(G2337GAT_737_gat) );
AND2XL U_g707 (.A(G2277GAT_714_ngat), .B(G2230GAT_697_ngat), .Y(G2330GAT_738_gat) );
AND2XL U_g708 (.A(G2171GAT_671_ngat), .B(G2285GAT_712_ngat), .Y(G2335GAT_739_gat) );
AND2XL U_g709 (.A(G2273GAT_715_ngat), .B(G2227GAT_698_ngat), .Y(G2328GAT_740_gat) );
AND2XL U_g710 (.A(G2166GAT_674_ngat), .B(G2281GAT_713_ngat), .Y(G2333GAT_741_gat) );
AND2XL U_g711 (.A(G2269GAT_716_ngat), .B(G2224GAT_699_ngat), .Y(G2326GAT_742_gat) );
AND2XL U_g712 (.A(G2161GAT_677_ngat), .B(G2277GAT_714_ngat), .Y(G2331GAT_743_gat) );
AND2XL U_g713 (.A(G2156GAT_680_ngat), .B(G2273GAT_715_ngat), .Y(G2329GAT_744_gat) );
AND2XL U_g714 (.A(G2151GAT_682_ngat), .B(G2269GAT_716_ngat), .Y(G2327GAT_745_gat) );
AND2XL U_g715 (.A(G2359GAT_717_ngat), .B(G1275GAT_43_ngat), .Y(G2410GAT_746_gat) );
AND2XL U_g716 (.A(G2358GAT_721_ngat), .B(G2357GAT_718_ngat), .Y(G2407GAT_747_gat) );
AND2XL U_g717 (.A(G2353GAT_723_ngat), .B(G2217GAT_643_ngat), .Y(G2404GAT_748_gat) );
AND2XL U_g718 (.A(G2353GAT_723_ngat), .B(G2319GAT_701_ngat), .Y(G2402GAT_749_gat) );
AND2XL U_g719 (.A(G2349GAT_725_ngat), .B(G2348GAT_720_ngat), .Y(G2395GAT_750_gat) );
AND2XL U_g720 (.A(G2347GAT_727_ngat), .B(G2346GAT_722_ngat), .Y(G2392GAT_751_gat) );
AND2XL U_g721 (.A(G1179GAT_75_ngat), .B(G2353GAT_723_ngat), .Y(G2403GAT_752_gat) );
AND2XL U_g722 (.A(G2345GAT_729_ngat), .B(G2344GAT_724_ngat), .Y(G2389GAT_753_gat) );
AND2XL U_g723 (.A(G1131GAT_91_ngat), .B(G2350GAT_719_ngat), .Y(G2398GAT_754_gat) );
AND2XL U_g724 (.A(G2343GAT_731_ngat), .B(G2342GAT_726_ngat), .Y(G2386GAT_755_gat) );
AND2XL U_g725 (.A(G2341GAT_733_ngat), .B(G2340GAT_728_ngat), .Y(G2383GAT_756_gat) );
AND2XL U_g726 (.A(G2339GAT_735_ngat), .B(G2338GAT_730_ngat), .Y(G2380GAT_757_gat) );
AND2XL U_g727 (.A(G2337GAT_737_ngat), .B(G2336GAT_732_ngat), .Y(G2377GAT_758_gat) );
AND2XL U_g728 (.A(G2335GAT_739_ngat), .B(G2334GAT_734_ngat), .Y(G2374GAT_759_gat) );
AND2XL U_g729 (.A(G2333GAT_741_ngat), .B(G2332GAT_736_ngat), .Y(G2371GAT_760_gat) );
AND2XL U_g730 (.A(G2331GAT_743_ngat), .B(G2330GAT_738_ngat), .Y(G2368GAT_761_gat) );
AND2XL U_g731 (.A(G2329GAT_744_ngat), .B(G2328GAT_740_ngat), .Y(G2365GAT_762_gat) );
AND2XL U_g732 (.A(G2327GAT_745_ngat), .B(G2326GAT_742_ngat), .Y(G2362GAT_763_gat) );
AND2XL U_g733 (.A(G2410GAT_746_ngat), .B(G1275GAT_43_ngat), .Y(G2474GAT_764_gat) );
AND2XL U_g734 (.A(G2359GAT_717_ngat), .B(G2410GAT_746_ngat), .Y(G2475GAT_765_gat) );
AND2XL U_g735 (.A(G2404GAT_748_ngat), .B(G2407GAT_747_ngat), .Y(G2470GAT_766_gat) );
AND2XL U_g736 (.A(G2403GAT_752_ngat), .B(G2402GAT_749_ngat), .Y(G2467GAT_767_gat) );
AND2XL U_g737 (.A(G2398GAT_754_ngat), .B(G2260GAT_687_ngat), .Y(G2464GAT_768_gat) );
AND2XL U_g738 (.A(G2398GAT_754_ngat), .B(G2350GAT_719_ngat), .Y(G2462GAT_769_gat) );
AND2XL U_g739 (.A(G1131GAT_91_ngat), .B(G2398GAT_754_ngat), .Y(G2463GAT_770_gat) );
AND2XL U_g740 (.A(G1083GAT_107_ngat), .B(G2395GAT_750_ngat), .Y(G2458GAT_771_gat) );
AND2XL U_g741 (.A(G1035GAT_123_ngat), .B(G2392GAT_751_ngat), .Y(G2454GAT_772_gat) );
AND2XL U_g742 (.A(G987GAT_139_ngat), .B(G2389GAT_753_ngat), .Y(G2450GAT_773_gat) );
AND2XL U_g743 (.A(G939GAT_155_ngat), .B(G2386GAT_755_ngat), .Y(G2446GAT_774_gat) );
AND2XL U_g744 (.A(G891GAT_171_ngat), .B(G2383GAT_756_ngat), .Y(G2442GAT_775_gat) );
AND2XL U_g745 (.A(G843GAT_187_ngat), .B(G2380GAT_757_ngat), .Y(G2438GAT_776_gat) );
AND2XL U_g746 (.A(G795GAT_203_ngat), .B(G2377GAT_758_ngat), .Y(G2434GAT_777_gat) );
AND2XL U_g747 (.A(G747GAT_219_ngat), .B(G2374GAT_759_ngat), .Y(G2430GAT_778_gat) );
AND2XL U_g748 (.A(G699GAT_235_ngat), .B(G2371GAT_760_ngat), .Y(G2426GAT_779_gat) );
AND2XL U_g749 (.A(G651GAT_251_ngat), .B(G2368GAT_761_ngat), .Y(G2422GAT_780_gat) );
AND2XL U_g750 (.A(G603GAT_267_ngat), .B(G2365GAT_762_ngat), .Y(G2418GAT_781_gat) );
AND2XL U_g751 (.A(G555GAT_283_ngat), .B(G2362GAT_763_ngat), .Y(G2414GAT_782_gat) );
AND2XL U_g752 (.A(G2475GAT_765_ngat), .B(G2474GAT_764_ngat), .Y(G2545GAT_783_gat) );
AND2XL U_g753 (.A(G2470GAT_766_ngat), .B(G2407GAT_747_ngat), .Y(G2543GAT_784_gat) );
AND2XL U_g754 (.A(G2404GAT_748_ngat), .B(G2470GAT_766_ngat), .Y(G2544GAT_785_gat) );
AND2XL U_g755 (.A(G2464GAT_768_ngat), .B(G2467GAT_767_ngat), .Y(G2539GAT_786_gat) );
AND2XL U_g756 (.A(G2463GAT_770_ngat), .B(G2462GAT_769_ngat), .Y(G2536GAT_787_gat) );
AND2XL U_g757 (.A(G2458GAT_771_ngat), .B(G2395GAT_750_ngat), .Y(G2531GAT_788_gat) );
AND2XL U_g758 (.A(G2454GAT_772_ngat), .B(G2392GAT_751_ngat), .Y(G2526GAT_789_gat) );
AND2XL U_g759 (.A(G2450GAT_773_ngat), .B(G2389GAT_753_ngat), .Y(G2521GAT_790_gat) );
AND2XL U_g760 (.A(G2458GAT_771_ngat), .B(G2313GAT_705_ngat), .Y(G2533GAT_791_gat) );
AND2XL U_g761 (.A(G2446GAT_774_ngat), .B(G2386GAT_755_ngat), .Y(G2516GAT_792_gat) );
AND2XL U_g762 (.A(G1083GAT_107_ngat), .B(G2458GAT_771_ngat), .Y(G2532GAT_793_gat) );
AND2XL U_g763 (.A(G2454GAT_772_ngat), .B(G2309GAT_706_ngat), .Y(G2528GAT_794_gat) );
AND2XL U_g764 (.A(G2442GAT_775_ngat), .B(G2383GAT_756_ngat), .Y(G2511GAT_795_gat) );
AND2XL U_g765 (.A(G1035GAT_123_ngat), .B(G2454GAT_772_ngat), .Y(G2527GAT_796_gat) );
AND2XL U_g766 (.A(G2450GAT_773_ngat), .B(G2305GAT_707_ngat), .Y(G2523GAT_797_gat) );
AND2XL U_g767 (.A(G2438GAT_776_ngat), .B(G2380GAT_757_ngat), .Y(G2506GAT_798_gat) );
AND2XL U_g768 (.A(G987GAT_139_ngat), .B(G2450GAT_773_ngat), .Y(G2522GAT_799_gat) );
AND2XL U_g769 (.A(G2446GAT_774_ngat), .B(G2301GAT_708_ngat), .Y(G2518GAT_800_gat) );
AND2XL U_g770 (.A(G2434GAT_777_ngat), .B(G2377GAT_758_ngat), .Y(G2501GAT_801_gat) );
AND2XL U_g771 (.A(G939GAT_155_ngat), .B(G2446GAT_774_ngat), .Y(G2517GAT_802_gat) );
AND2XL U_g772 (.A(G2442GAT_775_ngat), .B(G2297GAT_709_ngat), .Y(G2513GAT_803_gat) );
AND2XL U_g773 (.A(G2430GAT_778_ngat), .B(G2374GAT_759_ngat), .Y(G2496GAT_804_gat) );
AND2XL U_g774 (.A(G891GAT_171_ngat), .B(G2442GAT_775_ngat), .Y(G2512GAT_805_gat) );
AND2XL U_g775 (.A(G2438GAT_776_ngat), .B(G2293GAT_710_ngat), .Y(G2508GAT_806_gat) );
AND2XL U_g776 (.A(G2426GAT_779_ngat), .B(G2371GAT_760_ngat), .Y(G2491GAT_807_gat) );
AND2XL U_g777 (.A(G843GAT_187_ngat), .B(G2438GAT_776_ngat), .Y(G2507GAT_808_gat) );
AND2XL U_g778 (.A(G2434GAT_777_ngat), .B(G2289GAT_711_ngat), .Y(G2503GAT_809_gat) );
AND2XL U_g779 (.A(G2422GAT_780_ngat), .B(G2368GAT_761_ngat), .Y(G2486GAT_810_gat) );
AND2XL U_g780 (.A(G795GAT_203_ngat), .B(G2434GAT_777_ngat), .Y(G2502GAT_811_gat) );
AND2XL U_g781 (.A(G2430GAT_778_ngat), .B(G2285GAT_712_ngat), .Y(G2498GAT_812_gat) );
AND2XL U_g782 (.A(G2418GAT_781_ngat), .B(G2365GAT_762_ngat), .Y(G2481GAT_813_gat) );
AND2XL U_g783 (.A(G747GAT_219_ngat), .B(G2430GAT_778_ngat), .Y(G2497GAT_814_gat) );
AND2XL U_g784 (.A(G2426GAT_779_ngat), .B(G2281GAT_713_ngat), .Y(G2493GAT_815_gat) );
AND2XL U_g785 (.A(G2414GAT_782_ngat), .B(G2362GAT_763_ngat), .Y(G2476GAT_816_gat) );
AND2XL U_g786 (.A(G699GAT_235_ngat), .B(G2426GAT_779_ngat), .Y(G2492GAT_817_gat) );
AND2XL U_g787 (.A(G2422GAT_780_ngat), .B(G2277GAT_714_ngat), .Y(G2488GAT_818_gat) );
AND2XL U_g788 (.A(G651GAT_251_ngat), .B(G2422GAT_780_ngat), .Y(G2487GAT_819_gat) );
AND2XL U_g789 (.A(G2418GAT_781_ngat), .B(G2273GAT_715_ngat), .Y(G2483GAT_820_gat) );
AND2XL U_g790 (.A(G603GAT_267_ngat), .B(G2418GAT_781_ngat), .Y(G2482GAT_821_gat) );
AND2XL U_g791 (.A(G2414GAT_782_ngat), .B(G2269GAT_716_ngat), .Y(G2478GAT_822_gat) );
AND2XL U_g792 (.A(G555GAT_283_ngat), .B(G2414GAT_782_ngat), .Y(G2477GAT_823_gat) );
AND2XL U_g793 (.A(G2544GAT_785_ngat), .B(G2543GAT_784_ngat), .Y(G2588GAT_824_gat) );
AND2XL U_g794 (.A(G2539GAT_786_ngat), .B(G2467GAT_767_ngat), .Y(G2586GAT_825_gat) );
AND2XL U_g795 (.A(G2464GAT_768_ngat), .B(G2539GAT_786_ngat), .Y(G2587GAT_826_gat) );
AND2XL U_g796 (.A(G2533GAT_791_ngat), .B(G2536GAT_787_ngat), .Y(G2582GAT_827_gat) );
AND2XL U_g797 (.A(G2532GAT_793_ngat), .B(G2531GAT_788_ngat), .Y(G2579GAT_828_gat) );
AND2XL U_g798 (.A(G1230GAT_58_ngat), .B(G2545GAT_783_ngat), .Y(G2591GAT_829_gat) );
AND2XL U_g799 (.A(G2527GAT_796_ngat), .B(G2526GAT_789_ngat), .Y(G2576GAT_830_gat) );
AND2XL U_g800 (.A(G2522GAT_799_ngat), .B(G2521GAT_790_ngat), .Y(G2573GAT_831_gat) );
AND2XL U_g801 (.A(G2517GAT_802_ngat), .B(G2516GAT_792_ngat), .Y(G2570GAT_832_gat) );
AND2XL U_g802 (.A(G2512GAT_805_ngat), .B(G2511GAT_795_ngat), .Y(G2567GAT_833_gat) );
AND2XL U_g803 (.A(G2507GAT_808_ngat), .B(G2506GAT_798_ngat), .Y(G2564GAT_834_gat) );
AND2XL U_g804 (.A(G2502GAT_811_ngat), .B(G2501GAT_801_ngat), .Y(G2561GAT_835_gat) );
AND2XL U_g805 (.A(G2497GAT_814_ngat), .B(G2496GAT_804_ngat), .Y(G2558GAT_836_gat) );
AND2XL U_g806 (.A(G2492GAT_817_ngat), .B(G2491GAT_807_ngat), .Y(G2555GAT_837_gat) );
AND2XL U_g807 (.A(G2487GAT_819_ngat), .B(G2486GAT_810_ngat), .Y(G2552GAT_838_gat) );
AND2XL U_g808 (.A(G2482GAT_821_ngat), .B(G2481GAT_813_ngat), .Y(G2549GAT_839_gat) );
AND2XL U_g809 (.A(G2477GAT_823_ngat), .B(G2476GAT_816_ngat), .Y(G2548GAT_840_gat) );
AND2XL U_g810 (.A(G2591GAT_829_ngat), .B(G2410GAT_746_ngat), .Y(G2650GAT_841_gat) );
AND2XL U_g811 (.A(G2591GAT_829_ngat), .B(G2545GAT_783_ngat), .Y(G2648GAT_842_gat) );
AND2XL U_g812 (.A(G2587GAT_826_ngat), .B(G2586GAT_825_ngat), .Y(G2641GAT_843_gat) );
AND2XL U_g813 (.A(G2582GAT_827_ngat), .B(G2536GAT_787_ngat), .Y(G2639GAT_844_gat) );
AND2XL U_g814 (.A(G1230GAT_58_ngat), .B(G2591GAT_829_ngat), .Y(G2649GAT_845_gat) );
AND2XL U_g815 (.A(G1182GAT_74_ngat), .B(G2588GAT_824_ngat), .Y(G2644GAT_846_gat) );
AND2XL U_g816 (.A(G2533GAT_791_ngat), .B(G2582GAT_827_ngat), .Y(G2640GAT_847_gat) );
AND2XL U_g817 (.A(G2528GAT_794_ngat), .B(G2579GAT_828_ngat), .Y(G2635GAT_848_gat) );
AND2XL U_g818 (.A(G2523GAT_797_ngat), .B(G2576GAT_830_ngat), .Y(G2631GAT_849_gat) );
AND2XL U_g819 (.A(G2518GAT_800_ngat), .B(G2573GAT_831_ngat), .Y(G2627GAT_850_gat) );
AND2XL U_g820 (.A(G2513GAT_803_ngat), .B(G2570GAT_832_ngat), .Y(G2623GAT_851_gat) );
AND2XL U_g821 (.A(G2508GAT_806_ngat), .B(G2567GAT_833_ngat), .Y(G2619GAT_852_gat) );
AND2XL U_g822 (.A(G2503GAT_809_ngat), .B(G2564GAT_834_ngat), .Y(G2615GAT_853_gat) );
AND2XL U_g823 (.A(G2498GAT_812_ngat), .B(G2561GAT_835_ngat), .Y(G2611GAT_854_gat) );
AND2XL U_g824 (.A(G2493GAT_815_ngat), .B(G2558GAT_836_ngat), .Y(G2607GAT_855_gat) );
AND2XL U_g825 (.A(G2488GAT_818_ngat), .B(G2555GAT_837_ngat), .Y(G2603GAT_856_gat) );
AND2XL U_g826 (.A(G2483GAT_820_ngat), .B(G2552GAT_838_ngat), .Y(G2599GAT_857_gat) );
AND2XL U_g827 (.A(G2478GAT_822_ngat), .B(G2549GAT_839_ngat), .Y(G2595GAT_858_gat) );
AND2XL U_g828 (.A(G2650GAT_841_ngat), .B(G1278GAT_42_ngat), .Y(G2690GAT_859_gat) );
AND2XL U_g829 (.A(G2649GAT_845_ngat), .B(G2648GAT_842_ngat), .Y(G2687GAT_860_gat) );
AND2XL U_g830 (.A(G2644GAT_846_ngat), .B(G2470GAT_766_ngat), .Y(G2684GAT_861_gat) );
AND2XL U_g831 (.A(G2644GAT_846_ngat), .B(G2588GAT_824_ngat), .Y(G2682GAT_862_gat) );
AND2XL U_g832 (.A(G2640GAT_847_ngat), .B(G2639GAT_844_ngat), .Y(G2675GAT_863_gat) );
AND2XL U_g833 (.A(G2635GAT_848_ngat), .B(G2579GAT_828_ngat), .Y(G2673GAT_864_gat) );
AND2XL U_g834 (.A(G2631GAT_849_ngat), .B(G2576GAT_830_ngat), .Y(G2671GAT_865_gat) );
AND2XL U_g835 (.A(G1182GAT_74_ngat), .B(G2644GAT_846_ngat), .Y(G2683GAT_866_gat) );
AND2XL U_g836 (.A(G2627GAT_850_ngat), .B(G2573GAT_831_ngat), .Y(G2669GAT_867_gat) );
AND2XL U_g837 (.A(G1134GAT_90_ngat), .B(G2641GAT_843_ngat), .Y(G2678GAT_868_gat) );
AND2XL U_g838 (.A(G2623GAT_851_ngat), .B(G2570GAT_832_ngat), .Y(G2667GAT_869_gat) );
AND2XL U_g839 (.A(G2528GAT_794_ngat), .B(G2635GAT_848_ngat), .Y(G2674GAT_870_gat) );
AND2XL U_g840 (.A(G2619GAT_852_ngat), .B(G2567GAT_833_ngat), .Y(G2665GAT_871_gat) );
AND2XL U_g841 (.A(G2523GAT_797_ngat), .B(G2631GAT_849_ngat), .Y(G2672GAT_872_gat) );
AND2XL U_g842 (.A(G2615GAT_853_ngat), .B(G2564GAT_834_ngat), .Y(G2663GAT_873_gat) );
AND2XL U_g843 (.A(G2518GAT_800_ngat), .B(G2627GAT_850_ngat), .Y(G2670GAT_874_gat) );
AND2XL U_g844 (.A(G2611GAT_854_ngat), .B(G2561GAT_835_ngat), .Y(G2661GAT_875_gat) );
AND2XL U_g845 (.A(G2513GAT_803_ngat), .B(G2623GAT_851_ngat), .Y(G2668GAT_876_gat) );
AND2XL U_g846 (.A(G2607GAT_855_ngat), .B(G2558GAT_836_ngat), .Y(G2659GAT_877_gat) );
AND2XL U_g847 (.A(G2508GAT_806_ngat), .B(G2619GAT_852_ngat), .Y(G2666GAT_878_gat) );
AND2XL U_g848 (.A(G2603GAT_856_ngat), .B(G2555GAT_837_ngat), .Y(G2657GAT_879_gat) );
AND2XL U_g849 (.A(G2503GAT_809_ngat), .B(G2615GAT_853_ngat), .Y(G2664GAT_880_gat) );
AND2XL U_g850 (.A(G2599GAT_857_ngat), .B(G2552GAT_838_ngat), .Y(G2655GAT_881_gat) );
AND2XL U_g851 (.A(G2498GAT_812_ngat), .B(G2611GAT_854_ngat), .Y(G2662GAT_882_gat) );
AND2XL U_g852 (.A(G2595GAT_858_ngat), .B(G2549GAT_839_ngat), .Y(G2653GAT_883_gat) );
AND2XL U_g853 (.A(G2493GAT_815_ngat), .B(G2607GAT_855_ngat), .Y(G2660GAT_884_gat) );
AND2XL U_g854 (.A(G2488GAT_818_ngat), .B(G2603GAT_856_ngat), .Y(G2658GAT_885_gat) );
AND2XL U_g855 (.A(G2483GAT_820_ngat), .B(G2599GAT_857_ngat), .Y(G2656GAT_886_gat) );
AND2XL U_g856 (.A(G2478GAT_822_ngat), .B(G2595GAT_858_ngat), .Y(G2654GAT_887_gat) );
AND2XL U_g857 (.A(G2690GAT_859_ngat), .B(G1278GAT_42_ngat), .Y(G2743GAT_888_gat) );
AND2XL U_g858 (.A(G2650GAT_841_ngat), .B(G2690GAT_859_ngat), .Y(G2744GAT_889_gat) );
AND2XL U_g859 (.A(G2684GAT_861_ngat), .B(G2687GAT_860_ngat), .Y(G2739GAT_890_gat) );
AND2XL U_g860 (.A(G2683GAT_866_ngat), .B(G2682GAT_862_ngat), .Y(G2736GAT_891_gat) );
AND2XL U_g861 (.A(G2678GAT_868_ngat), .B(G2539GAT_786_ngat), .Y(G2733GAT_892_gat) );
AND2XL U_g862 (.A(G2678GAT_868_ngat), .B(G2641GAT_843_ngat), .Y(G2731GAT_893_gat) );
AND2XL U_g863 (.A(G2674GAT_870_ngat), .B(G2673GAT_864_ngat), .Y(G2724GAT_894_gat) );
AND2XL U_g864 (.A(G2672GAT_872_ngat), .B(G2671GAT_865_ngat), .Y(G2721GAT_895_gat) );
AND2XL U_g865 (.A(G2670GAT_874_ngat), .B(G2669GAT_867_ngat), .Y(G2718GAT_896_gat) );
AND2XL U_g866 (.A(G1134GAT_90_ngat), .B(G2678GAT_868_ngat), .Y(G2732GAT_897_gat) );
AND2XL U_g867 (.A(G2668GAT_876_ngat), .B(G2667GAT_869_ngat), .Y(G2715GAT_898_gat) );
AND2XL U_g868 (.A(G1086GAT_106_ngat), .B(G2675GAT_863_ngat), .Y(G2727GAT_899_gat) );
AND2XL U_g869 (.A(G2666GAT_878_ngat), .B(G2665GAT_871_ngat), .Y(G2712GAT_900_gat) );
AND2XL U_g870 (.A(G2664GAT_880_ngat), .B(G2663GAT_873_ngat), .Y(G2709GAT_901_gat) );
AND2XL U_g871 (.A(G2662GAT_882_ngat), .B(G2661GAT_875_ngat), .Y(G2706GAT_902_gat) );
AND2XL U_g872 (.A(G2660GAT_884_ngat), .B(G2659GAT_877_ngat), .Y(G2703GAT_903_gat) );
AND2XL U_g873 (.A(G2658GAT_885_ngat), .B(G2657GAT_879_ngat), .Y(G2700GAT_904_gat) );
AND2XL U_g874 (.A(G2656GAT_886_ngat), .B(G2655GAT_881_ngat), .Y(G2697GAT_905_gat) );
AND2XL U_g875 (.A(G2654GAT_887_ngat), .B(G2653GAT_883_ngat), .Y(G2694GAT_906_gat) );
AND2XL U_g876 (.A(G2744GAT_889_ngat), .B(G2743GAT_888_ngat), .Y(G2803GAT_907_gat) );
AND2XL U_g877 (.A(G2739GAT_890_ngat), .B(G2687GAT_860_ngat), .Y(G2801GAT_908_gat) );
AND2XL U_g878 (.A(G2684GAT_861_ngat), .B(G2739GAT_890_ngat), .Y(G2802GAT_909_gat) );
AND2XL U_g879 (.A(G2733GAT_892_ngat), .B(G2736GAT_891_ngat), .Y(G2797GAT_910_gat) );
AND2XL U_g880 (.A(G2732GAT_897_ngat), .B(G2731GAT_893_ngat), .Y(G2794GAT_911_gat) );
AND2XL U_g881 (.A(G2727GAT_899_ngat), .B(G2582GAT_827_ngat), .Y(G2791GAT_912_gat) );
AND2XL U_g882 (.A(G2727GAT_899_ngat), .B(G2675GAT_863_ngat), .Y(G2789GAT_913_gat) );
AND2XL U_g883 (.A(G1086GAT_106_ngat), .B(G2727GAT_899_ngat), .Y(G2790GAT_914_gat) );
AND2XL U_g884 (.A(G1038GAT_122_ngat), .B(G2724GAT_894_ngat), .Y(G2785GAT_915_gat) );
AND2XL U_g885 (.A(G990GAT_138_ngat), .B(G2721GAT_895_ngat), .Y(G2781GAT_916_gat) );
AND2XL U_g886 (.A(G942GAT_154_ngat), .B(G2718GAT_896_ngat), .Y(G2777GAT_917_gat) );
AND2XL U_g887 (.A(G894GAT_170_ngat), .B(G2715GAT_898_ngat), .Y(G2773GAT_918_gat) );
AND2XL U_g888 (.A(G846GAT_186_ngat), .B(G2712GAT_900_ngat), .Y(G2769GAT_919_gat) );
AND2XL U_g889 (.A(G798GAT_202_ngat), .B(G2709GAT_901_ngat), .Y(G2765GAT_920_gat) );
AND2XL U_g890 (.A(G750GAT_218_ngat), .B(G2706GAT_902_ngat), .Y(G2761GAT_921_gat) );
AND2XL U_g891 (.A(G702GAT_234_ngat), .B(G2703GAT_903_ngat), .Y(G2757GAT_922_gat) );
AND2XL U_g892 (.A(G654GAT_250_ngat), .B(G2700GAT_904_ngat), .Y(G2753GAT_923_gat) );
AND2XL U_g893 (.A(G606GAT_266_ngat), .B(G2697GAT_905_ngat), .Y(G2749GAT_924_gat) );
AND2XL U_g894 (.A(G558GAT_282_ngat), .B(G2694GAT_906_ngat), .Y(G2745GAT_925_gat) );
AND2XL U_g895 (.A(G2802GAT_909_ngat), .B(G2801GAT_908_ngat), .Y(G2870GAT_926_gat) );
AND2XL U_g896 (.A(G2797GAT_910_ngat), .B(G2736GAT_891_ngat), .Y(G2868GAT_927_gat) );
AND2XL U_g897 (.A(G2733GAT_892_ngat), .B(G2797GAT_910_ngat), .Y(G2869GAT_928_gat) );
AND2XL U_g898 (.A(G2791GAT_912_ngat), .B(G2794GAT_911_ngat), .Y(G2864GAT_929_gat) );
AND2XL U_g899 (.A(G2790GAT_914_ngat), .B(G2789GAT_913_ngat), .Y(G2861GAT_930_gat) );
AND2XL U_g900 (.A(G2785GAT_915_ngat), .B(G2724GAT_894_ngat), .Y(G2856GAT_931_gat) );
AND2XL U_g901 (.A(G1233GAT_57_ngat), .B(G2803GAT_907_ngat), .Y(G2873GAT_932_gat) );
AND2XL U_g902 (.A(G2781GAT_916_ngat), .B(G2721GAT_895_ngat), .Y(G2851GAT_933_gat) );
AND2XL U_g903 (.A(G2777GAT_917_ngat), .B(G2718GAT_896_ngat), .Y(G2846GAT_934_gat) );
AND2XL U_g904 (.A(G2773GAT_918_ngat), .B(G2715GAT_898_ngat), .Y(G2841GAT_935_gat) );
AND2XL U_g905 (.A(G2785GAT_915_ngat), .B(G2635GAT_848_ngat), .Y(G2858GAT_936_gat) );
AND2XL U_g906 (.A(G2769GAT_919_ngat), .B(G2712GAT_900_ngat), .Y(G2836GAT_937_gat) );
AND2XL U_g907 (.A(G1038GAT_122_ngat), .B(G2785GAT_915_ngat), .Y(G2857GAT_938_gat) );
AND2XL U_g908 (.A(G2781GAT_916_ngat), .B(G2631GAT_849_ngat), .Y(G2853GAT_939_gat) );
AND2XL U_g909 (.A(G2765GAT_920_ngat), .B(G2709GAT_901_ngat), .Y(G2831GAT_940_gat) );
AND2XL U_g910 (.A(G990GAT_138_ngat), .B(G2781GAT_916_ngat), .Y(G2852GAT_941_gat) );
AND2XL U_g911 (.A(G2777GAT_917_ngat), .B(G2627GAT_850_ngat), .Y(G2848GAT_942_gat) );
AND2XL U_g912 (.A(G2761GAT_921_ngat), .B(G2706GAT_902_ngat), .Y(G2826GAT_943_gat) );
AND2XL U_g913 (.A(G942GAT_154_ngat), .B(G2777GAT_917_ngat), .Y(G2847GAT_944_gat) );
AND2XL U_g914 (.A(G2773GAT_918_ngat), .B(G2623GAT_851_ngat), .Y(G2843GAT_945_gat) );
AND2XL U_g915 (.A(G2757GAT_922_ngat), .B(G2703GAT_903_ngat), .Y(G2821GAT_946_gat) );
AND2XL U_g916 (.A(G894GAT_170_ngat), .B(G2773GAT_918_ngat), .Y(G2842GAT_947_gat) );
AND2XL U_g917 (.A(G2769GAT_919_ngat), .B(G2619GAT_852_ngat), .Y(G2838GAT_948_gat) );
AND2XL U_g918 (.A(G2753GAT_923_ngat), .B(G2700GAT_904_ngat), .Y(G2816GAT_949_gat) );
AND2XL U_g919 (.A(G846GAT_186_ngat), .B(G2769GAT_919_ngat), .Y(G2837GAT_950_gat) );
AND2XL U_g920 (.A(G2765GAT_920_ngat), .B(G2615GAT_853_ngat), .Y(G2833GAT_951_gat) );
AND2XL U_g921 (.A(G2749GAT_924_ngat), .B(G2697GAT_905_ngat), .Y(G2811GAT_952_gat) );
AND2XL U_g922 (.A(G798GAT_202_ngat), .B(G2765GAT_920_ngat), .Y(G2832GAT_953_gat) );
AND2XL U_g923 (.A(G2761GAT_921_ngat), .B(G2611GAT_854_ngat), .Y(G2828GAT_954_gat) );
AND2XL U_g924 (.A(G2745GAT_925_ngat), .B(G2694GAT_906_ngat), .Y(G2806GAT_955_gat) );
AND2XL U_g925 (.A(G750GAT_218_ngat), .B(G2761GAT_921_ngat), .Y(G2827GAT_956_gat) );
AND2XL U_g926 (.A(G2757GAT_922_ngat), .B(G2607GAT_855_ngat), .Y(G2823GAT_957_gat) );
AND2XL U_g927 (.A(G702GAT_234_ngat), .B(G2757GAT_922_ngat), .Y(G2822GAT_958_gat) );
AND2XL U_g928 (.A(G2753GAT_923_ngat), .B(G2603GAT_856_ngat), .Y(G2818GAT_959_gat) );
AND2XL U_g929 (.A(G654GAT_250_ngat), .B(G2753GAT_923_ngat), .Y(G2817GAT_960_gat) );
AND2XL U_g930 (.A(G2749GAT_924_ngat), .B(G2599GAT_857_ngat), .Y(G2813GAT_961_gat) );
AND2XL U_g931 (.A(G606GAT_266_ngat), .B(G2749GAT_924_ngat), .Y(G2812GAT_962_gat) );
AND2XL U_g932 (.A(G2745GAT_925_ngat), .B(G2595GAT_858_ngat), .Y(G2808GAT_963_gat) );
AND2XL U_g933 (.A(G558GAT_282_ngat), .B(G2745GAT_925_ngat), .Y(G2807GAT_964_gat) );
AND2XL U_g934 (.A(G2873GAT_932_ngat), .B(G2690GAT_859_ngat), .Y(G2923GAT_965_gat) );
AND2XL U_g935 (.A(G2873GAT_932_ngat), .B(G2803GAT_907_ngat), .Y(G2921GAT_966_gat) );
AND2XL U_g936 (.A(G2869GAT_928_ngat), .B(G2868GAT_927_ngat), .Y(G2914GAT_967_gat) );
AND2XL U_g937 (.A(G2864GAT_929_ngat), .B(G2794GAT_911_ngat), .Y(G2912GAT_968_gat) );
AND2XL U_g938 (.A(G2791GAT_912_ngat), .B(G2864GAT_929_ngat), .Y(G2913GAT_969_gat) );
AND2XL U_g939 (.A(G2858GAT_936_ngat), .B(G2861GAT_930_ngat), .Y(G2908GAT_970_gat) );
AND2XL U_g940 (.A(G2857GAT_938_ngat), .B(G2856GAT_931_ngat), .Y(G2905GAT_971_gat) );
AND2XL U_g941 (.A(G1233GAT_57_ngat), .B(G2873GAT_932_ngat), .Y(G2922GAT_972_gat) );
AND2XL U_g942 (.A(G2852GAT_941_ngat), .B(G2851GAT_933_ngat), .Y(G2902GAT_973_gat) );
AND2XL U_g943 (.A(G1185GAT_73_ngat), .B(G2870GAT_926_ngat), .Y(G2917GAT_974_gat) );
AND2XL U_g944 (.A(G2847GAT_944_ngat), .B(G2846GAT_934_ngat), .Y(G2899GAT_975_gat) );
AND2XL U_g945 (.A(G2842GAT_947_ngat), .B(G2841GAT_935_ngat), .Y(G2896GAT_976_gat) );
AND2XL U_g946 (.A(G2837GAT_950_ngat), .B(G2836GAT_937_ngat), .Y(G2893GAT_977_gat) );
AND2XL U_g947 (.A(G2832GAT_953_ngat), .B(G2831GAT_940_ngat), .Y(G2890GAT_978_gat) );
AND2XL U_g948 (.A(G2827GAT_956_ngat), .B(G2826GAT_943_ngat), .Y(G2887GAT_979_gat) );
AND2XL U_g949 (.A(G2822GAT_958_ngat), .B(G2821GAT_946_ngat), .Y(G2884GAT_980_gat) );
AND2XL U_g950 (.A(G2817GAT_960_ngat), .B(G2816GAT_949_ngat), .Y(G2881GAT_981_gat) );
AND2XL U_g951 (.A(G2812GAT_962_ngat), .B(G2811GAT_952_ngat), .Y(G2878GAT_982_gat) );
AND2XL U_g952 (.A(G2807GAT_964_ngat), .B(G2806GAT_955_ngat), .Y(G2877GAT_983_gat) );
AND2XL U_g953 (.A(G2923GAT_965_ngat), .B(G1281GAT_41_ngat), .Y(G2983GAT_984_gat) );
AND2XL U_g954 (.A(G2922GAT_972_ngat), .B(G2921GAT_966_ngat), .Y(G2980GAT_985_gat) );
AND2XL U_g955 (.A(G2917GAT_974_ngat), .B(G2739GAT_890_ngat), .Y(G2977GAT_986_gat) );
AND2XL U_g956 (.A(G2917GAT_974_ngat), .B(G2870GAT_926_ngat), .Y(G2975GAT_987_gat) );
AND2XL U_g957 (.A(G2913GAT_969_ngat), .B(G2912GAT_968_ngat), .Y(G2968GAT_988_gat) );
AND2XL U_g958 (.A(G2908GAT_970_ngat), .B(G2861GAT_930_ngat), .Y(G2966GAT_989_gat) );
AND2XL U_g959 (.A(G1185GAT_73_ngat), .B(G2917GAT_974_ngat), .Y(G2976GAT_990_gat) );
AND2XL U_g960 (.A(G1137GAT_89_ngat), .B(G2914GAT_967_ngat), .Y(G2971GAT_991_gat) );
AND2XL U_g961 (.A(G2858GAT_936_ngat), .B(G2908GAT_970_ngat), .Y(G2967GAT_992_gat) );
AND2XL U_g962 (.A(G2853GAT_939_ngat), .B(G2905GAT_971_ngat), .Y(G2962GAT_993_gat) );
AND2XL U_g963 (.A(G2848GAT_942_ngat), .B(G2902GAT_973_ngat), .Y(G2958GAT_994_gat) );
AND2XL U_g964 (.A(G2843GAT_945_ngat), .B(G2899GAT_975_ngat), .Y(G2954GAT_995_gat) );
AND2XL U_g965 (.A(G2838GAT_948_ngat), .B(G2896GAT_976_ngat), .Y(G2950GAT_996_gat) );
AND2XL U_g966 (.A(G2833GAT_951_ngat), .B(G2893GAT_977_ngat), .Y(G2946GAT_997_gat) );
AND2XL U_g967 (.A(G2828GAT_954_ngat), .B(G2890GAT_978_ngat), .Y(G2942GAT_998_gat) );
AND2XL U_g968 (.A(G2823GAT_957_ngat), .B(G2887GAT_979_ngat), .Y(G2938GAT_999_gat) );
AND2XL U_g969 (.A(G2818GAT_959_ngat), .B(G2884GAT_980_ngat), .Y(G2934GAT_1000_gat) );
AND2XL U_g970 (.A(G2813GAT_961_ngat), .B(G2881GAT_981_ngat), .Y(G2930GAT_1001_gat) );
AND2XL U_g971 (.A(G2808GAT_963_ngat), .B(G2878GAT_982_ngat), .Y(G2926GAT_1002_gat) );
AND2XL U_g972 (.A(G2983GAT_984_ngat), .B(G1281GAT_41_ngat), .Y(G3026GAT_1003_gat) );
AND2XL U_g973 (.A(G2923GAT_965_ngat), .B(G2983GAT_984_ngat), .Y(G3027GAT_1004_gat) );
AND2XL U_g974 (.A(G2977GAT_986_ngat), .B(G2980GAT_985_ngat), .Y(G3022GAT_1005_gat) );
AND2XL U_g975 (.A(G2976GAT_990_ngat), .B(G2975GAT_987_ngat), .Y(G3019GAT_1006_gat) );
AND2XL U_g976 (.A(G2971GAT_991_ngat), .B(G2797GAT_910_ngat), .Y(G3016GAT_1007_gat) );
AND2XL U_g977 (.A(G2971GAT_991_ngat), .B(G2914GAT_967_ngat), .Y(G3014GAT_1008_gat) );
AND2XL U_g978 (.A(G2967GAT_992_ngat), .B(G2966GAT_989_ngat), .Y(G3007GAT_1009_gat) );
AND2XL U_g979 (.A(G2962GAT_993_ngat), .B(G2905GAT_971_ngat), .Y(G3005GAT_1010_gat) );
AND2XL U_g980 (.A(G2958GAT_994_ngat), .B(G2902GAT_973_ngat), .Y(G3003GAT_1011_gat) );
AND2XL U_g981 (.A(G2954GAT_995_ngat), .B(G2899GAT_975_ngat), .Y(G3001GAT_1012_gat) );
AND2XL U_g982 (.A(G1137GAT_89_ngat), .B(G2971GAT_991_ngat), .Y(G3015GAT_1013_gat) );
AND2XL U_g983 (.A(G2950GAT_996_ngat), .B(G2896GAT_976_ngat), .Y(G2999GAT_1014_gat) );
AND2XL U_g984 (.A(G1089GAT_105_ngat), .B(G2968GAT_988_ngat), .Y(G3010GAT_1015_gat) );
AND2XL U_g985 (.A(G2946GAT_997_ngat), .B(G2893GAT_977_ngat), .Y(G2997GAT_1016_gat) );
AND2XL U_g986 (.A(G2853GAT_939_ngat), .B(G2962GAT_993_ngat), .Y(G3006GAT_1017_gat) );
AND2XL U_g987 (.A(G2942GAT_998_ngat), .B(G2890GAT_978_ngat), .Y(G2995GAT_1018_gat) );
AND2XL U_g988 (.A(G2848GAT_942_ngat), .B(G2958GAT_994_ngat), .Y(G3004GAT_1019_gat) );
AND2XL U_g989 (.A(G2938GAT_999_ngat), .B(G2887GAT_979_ngat), .Y(G2993GAT_1020_gat) );
AND2XL U_g990 (.A(G2843GAT_945_ngat), .B(G2954GAT_995_ngat), .Y(G3002GAT_1021_gat) );
AND2XL U_g991 (.A(G2934GAT_1000_ngat), .B(G2884GAT_980_ngat), .Y(G2991GAT_1022_gat) );
AND2XL U_g992 (.A(G2838GAT_948_ngat), .B(G2950GAT_996_ngat), .Y(G3000GAT_1023_gat) );
AND2XL U_g993 (.A(G2930GAT_1001_ngat), .B(G2881GAT_981_ngat), .Y(G2989GAT_1024_gat) );
AND2XL U_g994 (.A(G2833GAT_951_ngat), .B(G2946GAT_997_ngat), .Y(G2998GAT_1025_gat) );
AND2XL U_g995 (.A(G2926GAT_1002_ngat), .B(G2878GAT_982_ngat), .Y(G2987GAT_1026_gat) );
AND2XL U_g996 (.A(G2828GAT_954_ngat), .B(G2942GAT_998_ngat), .Y(G2996GAT_1027_gat) );
AND2XL U_g997 (.A(G2823GAT_957_ngat), .B(G2938GAT_999_ngat), .Y(G2994GAT_1028_gat) );
AND2XL U_g998 (.A(G2818GAT_959_ngat), .B(G2934GAT_1000_ngat), .Y(G2992GAT_1029_gat) );
AND2XL U_g999 (.A(G2813GAT_961_ngat), .B(G2930GAT_1001_ngat), .Y(G2990GAT_1030_gat) );
AND2XL U_g1000 (.A(G2808GAT_963_ngat), .B(G2926GAT_1002_ngat), .Y(G2988GAT_1031_gat) );
AND2XL U_g1001 (.A(G3027GAT_1004_ngat), .B(G3026GAT_1003_ngat), .Y(G3076GAT_1032_gat) );
AND2XL U_g1002 (.A(G3022GAT_1005_ngat), .B(G2980GAT_985_ngat), .Y(G3074GAT_1033_gat) );
AND2XL U_g1003 (.A(G2977GAT_986_ngat), .B(G3022GAT_1005_ngat), .Y(G3075GAT_1034_gat) );
AND2XL U_g1004 (.A(G3016GAT_1007_ngat), .B(G3019GAT_1006_ngat), .Y(G3070GAT_1035_gat) );
AND2XL U_g1005 (.A(G3015GAT_1013_ngat), .B(G3014GAT_1008_ngat), .Y(G3067GAT_1036_gat) );
AND2XL U_g1006 (.A(G3010GAT_1015_ngat), .B(G2864GAT_929_ngat), .Y(G3064GAT_1037_gat) );
AND2XL U_g1007 (.A(G3010GAT_1015_ngat), .B(G2968GAT_988_ngat), .Y(G3062GAT_1038_gat) );
AND2XL U_g1008 (.A(G3006GAT_1017_ngat), .B(G3005GAT_1010_ngat), .Y(G3055GAT_1039_gat) );
AND2XL U_g1009 (.A(G3004GAT_1019_ngat), .B(G3003GAT_1011_ngat), .Y(G3052GAT_1040_gat) );
AND2XL U_g1010 (.A(G3002GAT_1021_ngat), .B(G3001GAT_1012_ngat), .Y(G3049GAT_1041_gat) );
AND2XL U_g1011 (.A(G3000GAT_1023_ngat), .B(G2999GAT_1014_ngat), .Y(G3046GAT_1042_gat) );
AND2XL U_g1012 (.A(G1089GAT_105_ngat), .B(G3010GAT_1015_ngat), .Y(G3063GAT_1043_gat) );
AND2XL U_g1013 (.A(G2998GAT_1025_ngat), .B(G2997GAT_1016_ngat), .Y(G3043GAT_1044_gat) );
AND2XL U_g1014 (.A(G1041GAT_121_ngat), .B(G3007GAT_1009_ngat), .Y(G3058GAT_1045_gat) );
AND2XL U_g1015 (.A(G2996GAT_1027_ngat), .B(G2995GAT_1018_ngat), .Y(G3040GAT_1046_gat) );
AND2XL U_g1016 (.A(G2994GAT_1028_ngat), .B(G2993GAT_1020_ngat), .Y(G3037GAT_1047_gat) );
AND2XL U_g1017 (.A(G2992GAT_1029_ngat), .B(G2991GAT_1022_ngat), .Y(G3034GAT_1048_gat) );
AND2XL U_g1018 (.A(G2990GAT_1030_ngat), .B(G2989GAT_1024_ngat), .Y(G3031GAT_1049_gat) );
AND2XL U_g1019 (.A(G2988GAT_1031_ngat), .B(G2987GAT_1026_ngat), .Y(G3028GAT_1050_gat) );
AND2XL U_g1020 (.A(G3075GAT_1034_ngat), .B(G3074GAT_1033_ngat), .Y(G3133GAT_1051_gat) );
AND2XL U_g1021 (.A(G3070GAT_1035_ngat), .B(G3019GAT_1006_ngat), .Y(G3131GAT_1052_gat) );
AND2XL U_g1022 (.A(G3016GAT_1007_ngat), .B(G3070GAT_1035_ngat), .Y(G3132GAT_1053_gat) );
AND2XL U_g1023 (.A(G3064GAT_1037_ngat), .B(G3067GAT_1036_ngat), .Y(G3127GAT_1054_gat) );
AND2XL U_g1024 (.A(G3063GAT_1043_ngat), .B(G3062GAT_1038_ngat), .Y(G3124GAT_1055_gat) );
AND2XL U_g1025 (.A(G3058GAT_1045_ngat), .B(G2908GAT_970_ngat), .Y(G3121GAT_1056_gat) );
AND2XL U_g1026 (.A(G3058GAT_1045_ngat), .B(G3007GAT_1009_ngat), .Y(G3119GAT_1057_gat) );
AND2XL U_g1027 (.A(G1236GAT_56_ngat), .B(G3076GAT_1032_ngat), .Y(G3136GAT_1058_gat) );
AND2XL U_g1028 (.A(G1041GAT_121_ngat), .B(G3058GAT_1045_ngat), .Y(G3120GAT_1059_gat) );
AND2XL U_g1029 (.A(G993GAT_137_ngat), .B(G3055GAT_1039_ngat), .Y(G3115GAT_1060_gat) );
AND2XL U_g1030 (.A(G945GAT_153_ngat), .B(G3052GAT_1040_ngat), .Y(G3111GAT_1061_gat) );
AND2XL U_g1031 (.A(G897GAT_169_ngat), .B(G3049GAT_1041_ngat), .Y(G3107GAT_1062_gat) );
AND2XL U_g1032 (.A(G849GAT_185_ngat), .B(G3046GAT_1042_ngat), .Y(G3103GAT_1063_gat) );
AND2XL U_g1033 (.A(G801GAT_201_ngat), .B(G3043GAT_1044_ngat), .Y(G3099GAT_1064_gat) );
AND2XL U_g1034 (.A(G753GAT_217_ngat), .B(G3040GAT_1046_ngat), .Y(G3095GAT_1065_gat) );
AND2XL U_g1035 (.A(G705GAT_233_ngat), .B(G3037GAT_1047_ngat), .Y(G3091GAT_1066_gat) );
AND2XL U_g1036 (.A(G657GAT_249_ngat), .B(G3034GAT_1048_ngat), .Y(G3087GAT_1067_gat) );
AND2XL U_g1037 (.A(G609GAT_265_ngat), .B(G3031GAT_1049_ngat), .Y(G3083GAT_1068_gat) );
AND2XL U_g1038 (.A(G561GAT_281_ngat), .B(G3028GAT_1050_ngat), .Y(G3079GAT_1069_gat) );
AND2XL U_g1039 (.A(G3136GAT_1058_ngat), .B(G2983GAT_984_ngat), .Y(G3208GAT_1070_gat) );
AND2XL U_g1040 (.A(G3136GAT_1058_ngat), .B(G3076GAT_1032_ngat), .Y(G3206GAT_1071_gat) );
AND2XL U_g1041 (.A(G3132GAT_1053_ngat), .B(G3131GAT_1052_ngat), .Y(G3199GAT_1072_gat) );
AND2XL U_g1042 (.A(G3127GAT_1054_ngat), .B(G3067GAT_1036_ngat), .Y(G3197GAT_1073_gat) );
AND2XL U_g1043 (.A(G3064GAT_1037_ngat), .B(G3127GAT_1054_ngat), .Y(G3198GAT_1074_gat) );
AND2XL U_g1044 (.A(G3121GAT_1056_ngat), .B(G3124GAT_1055_ngat), .Y(G3193GAT_1075_gat) );
AND2XL U_g1045 (.A(G3120GAT_1059_ngat), .B(G3119GAT_1057_ngat), .Y(G3190GAT_1076_gat) );
AND2XL U_g1046 (.A(G3115GAT_1060_ngat), .B(G3055GAT_1039_ngat), .Y(G3185GAT_1077_gat) );
AND2XL U_g1047 (.A(G1236GAT_56_ngat), .B(G3136GAT_1058_ngat), .Y(G3207GAT_1078_gat) );
AND2XL U_g1048 (.A(G3111GAT_1061_ngat), .B(G3052GAT_1040_ngat), .Y(G3180GAT_1079_gat) );
AND2XL U_g1049 (.A(G1188GAT_72_ngat), .B(G3133GAT_1051_ngat), .Y(G3202GAT_1080_gat) );
AND2XL U_g1050 (.A(G3107GAT_1062_ngat), .B(G3049GAT_1041_ngat), .Y(G3175GAT_1081_gat) );
AND2XL U_g1051 (.A(G3103GAT_1063_ngat), .B(G3046GAT_1042_ngat), .Y(G3170GAT_1082_gat) );
AND2XL U_g1052 (.A(G3099GAT_1064_ngat), .B(G3043GAT_1044_ngat), .Y(G3165GAT_1083_gat) );
AND2XL U_g1053 (.A(G3115GAT_1060_ngat), .B(G2962GAT_993_ngat), .Y(G3187GAT_1084_gat) );
AND2XL U_g1054 (.A(G3095GAT_1065_ngat), .B(G3040GAT_1046_ngat), .Y(G3160GAT_1085_gat) );
AND2XL U_g1055 (.A(G993GAT_137_ngat), .B(G3115GAT_1060_ngat), .Y(G3186GAT_1086_gat) );
AND2XL U_g1056 (.A(G3111GAT_1061_ngat), .B(G2958GAT_994_ngat), .Y(G3182GAT_1087_gat) );
AND2XL U_g1057 (.A(G3091GAT_1066_ngat), .B(G3037GAT_1047_ngat), .Y(G3155GAT_1088_gat) );
AND2XL U_g1058 (.A(G945GAT_153_ngat), .B(G3111GAT_1061_ngat), .Y(G3181GAT_1089_gat) );
AND2XL U_g1059 (.A(G3107GAT_1062_ngat), .B(G2954GAT_995_ngat), .Y(G3177GAT_1090_gat) );
AND2XL U_g1060 (.A(G3087GAT_1067_ngat), .B(G3034GAT_1048_ngat), .Y(G3150GAT_1091_gat) );
AND2XL U_g1061 (.A(G897GAT_169_ngat), .B(G3107GAT_1062_ngat), .Y(G3176GAT_1092_gat) );
AND2XL U_g1062 (.A(G3103GAT_1063_ngat), .B(G2950GAT_996_ngat), .Y(G3172GAT_1093_gat) );
AND2XL U_g1063 (.A(G3083GAT_1068_ngat), .B(G3031GAT_1049_ngat), .Y(G3145GAT_1094_gat) );
AND2XL U_g1064 (.A(G849GAT_185_ngat), .B(G3103GAT_1063_ngat), .Y(G3171GAT_1095_gat) );
AND2XL U_g1065 (.A(G3099GAT_1064_ngat), .B(G2946GAT_997_ngat), .Y(G3167GAT_1096_gat) );
AND2XL U_g1066 (.A(G3079GAT_1069_ngat), .B(G3028GAT_1050_ngat), .Y(G3140GAT_1097_gat) );
AND2XL U_g1067 (.A(G801GAT_201_ngat), .B(G3099GAT_1064_ngat), .Y(G3166GAT_1098_gat) );
AND2XL U_g1068 (.A(G3095GAT_1065_ngat), .B(G2942GAT_998_ngat), .Y(G3162GAT_1099_gat) );
AND2XL U_g1069 (.A(G753GAT_217_ngat), .B(G3095GAT_1065_ngat), .Y(G3161GAT_1100_gat) );
AND2XL U_g1070 (.A(G3091GAT_1066_ngat), .B(G2938GAT_999_ngat), .Y(G3157GAT_1101_gat) );
AND2XL U_g1071 (.A(G705GAT_233_ngat), .B(G3091GAT_1066_ngat), .Y(G3156GAT_1102_gat) );
AND2XL U_g1072 (.A(G3087GAT_1067_ngat), .B(G2934GAT_1000_ngat), .Y(G3152GAT_1103_gat) );
AND2XL U_g1073 (.A(G657GAT_249_ngat), .B(G3087GAT_1067_ngat), .Y(G3151GAT_1104_gat) );
AND2XL U_g1074 (.A(G3083GAT_1068_ngat), .B(G2930GAT_1001_ngat), .Y(G3147GAT_1105_gat) );
AND2XL U_g1075 (.A(G609GAT_265_ngat), .B(G3083GAT_1068_ngat), .Y(G3146GAT_1106_gat) );
AND2XL U_g1076 (.A(G3079GAT_1069_ngat), .B(G2926GAT_1002_ngat), .Y(G3142GAT_1107_gat) );
AND2XL U_g1077 (.A(G561GAT_281_ngat), .B(G3079GAT_1069_ngat), .Y(G3141GAT_1108_gat) );
AND2XL U_g1078 (.A(G3208GAT_1070_ngat), .B(G1284GAT_40_ngat), .Y(G3260GAT_1109_gat) );
AND2XL U_g1079 (.A(G3207GAT_1078_ngat), .B(G3206GAT_1071_ngat), .Y(G3257GAT_1110_gat) );
AND2XL U_g1080 (.A(G3202GAT_1080_ngat), .B(G3022GAT_1005_ngat), .Y(G3254GAT_1111_gat) );
AND2XL U_g1081 (.A(G3202GAT_1080_ngat), .B(G3133GAT_1051_ngat), .Y(G3252GAT_1112_gat) );
AND2XL U_g1082 (.A(G3198GAT_1074_ngat), .B(G3197GAT_1073_ngat), .Y(G3245GAT_1113_gat) );
AND2XL U_g1083 (.A(G3193GAT_1075_ngat), .B(G3124GAT_1055_ngat), .Y(G3243GAT_1114_gat) );
AND2XL U_g1084 (.A(G3121GAT_1056_ngat), .B(G3193GAT_1075_ngat), .Y(G3244GAT_1115_gat) );
AND2XL U_g1085 (.A(G3187GAT_1084_ngat), .B(G3190GAT_1076_ngat), .Y(G3239GAT_1116_gat) );
AND2XL U_g1086 (.A(G3186GAT_1086_ngat), .B(G3185GAT_1077_ngat), .Y(G3236GAT_1117_gat) );
AND2XL U_g1087 (.A(G3181GAT_1089_ngat), .B(G3180GAT_1079_ngat), .Y(G3233GAT_1118_gat) );
AND2XL U_g1088 (.A(G1188GAT_72_ngat), .B(G3202GAT_1080_ngat), .Y(G3253GAT_1119_gat) );
AND2XL U_g1089 (.A(G3176GAT_1092_ngat), .B(G3175GAT_1081_ngat), .Y(G3230GAT_1120_gat) );
AND2XL U_g1090 (.A(G1140GAT_88_ngat), .B(G3199GAT_1072_ngat), .Y(G3248GAT_1121_gat) );
AND2XL U_g1091 (.A(G3171GAT_1095_ngat), .B(G3170GAT_1082_ngat), .Y(G3227GAT_1122_gat) );
AND2XL U_g1092 (.A(G3166GAT_1098_ngat), .B(G3165GAT_1083_ngat), .Y(G3224GAT_1123_gat) );
AND2XL U_g1093 (.A(G3161GAT_1100_ngat), .B(G3160GAT_1085_ngat), .Y(G3221GAT_1124_gat) );
AND2XL U_g1094 (.A(G3156GAT_1102_ngat), .B(G3155GAT_1088_ngat), .Y(G3218GAT_1125_gat) );
AND2XL U_g1095 (.A(G3151GAT_1104_ngat), .B(G3150GAT_1091_ngat), .Y(G3215GAT_1126_gat) );
AND2XL U_g1096 (.A(G3146GAT_1106_ngat), .B(G3145GAT_1094_ngat), .Y(G3212GAT_1127_gat) );
AND2XL U_g1097 (.A(G3141GAT_1108_ngat), .B(G3140GAT_1097_ngat), .Y(G3211GAT_1128_gat) );
AND2XL U_g1098 (.A(G3260GAT_1109_ngat), .B(G1284GAT_40_ngat), .Y(G3321GAT_1129_gat) );
AND2XL U_g1099 (.A(G3208GAT_1070_ngat), .B(G3260GAT_1109_ngat), .Y(G3322GAT_1130_gat) );
AND2XL U_g1100 (.A(G3254GAT_1111_ngat), .B(G3257GAT_1110_ngat), .Y(G3317GAT_1131_gat) );
AND2XL U_g1101 (.A(G3253GAT_1119_ngat), .B(G3252GAT_1112_ngat), .Y(G3314GAT_1132_gat) );
AND2XL U_g1102 (.A(G3248GAT_1121_ngat), .B(G3070GAT_1035_ngat), .Y(G3311GAT_1133_gat) );
AND2XL U_g1103 (.A(G3248GAT_1121_ngat), .B(G3199GAT_1072_ngat), .Y(G3309GAT_1134_gat) );
AND2XL U_g1104 (.A(G3244GAT_1115_ngat), .B(G3243GAT_1114_ngat), .Y(G3302GAT_1135_gat) );
AND2XL U_g1105 (.A(G3239GAT_1116_ngat), .B(G3190GAT_1076_ngat), .Y(G3300GAT_1136_gat) );
AND2XL U_g1106 (.A(G1140GAT_88_ngat), .B(G3248GAT_1121_ngat), .Y(G3310GAT_1137_gat) );
AND2XL U_g1107 (.A(G1092GAT_104_ngat), .B(G3245GAT_1113_ngat), .Y(G3305GAT_1138_gat) );
AND2XL U_g1108 (.A(G3187GAT_1084_ngat), .B(G3239GAT_1116_ngat), .Y(G3301GAT_1139_gat) );
AND2XL U_g1109 (.A(G3182GAT_1087_ngat), .B(G3236GAT_1117_ngat), .Y(G3296GAT_1140_gat) );
AND2XL U_g1110 (.A(G3177GAT_1090_ngat), .B(G3233GAT_1118_ngat), .Y(G3292GAT_1141_gat) );
AND2XL U_g1111 (.A(G3172GAT_1093_ngat), .B(G3230GAT_1120_ngat), .Y(G3288GAT_1142_gat) );
AND2XL U_g1112 (.A(G3167GAT_1096_ngat), .B(G3227GAT_1122_ngat), .Y(G3284GAT_1143_gat) );
AND2XL U_g1113 (.A(G3162GAT_1099_ngat), .B(G3224GAT_1123_ngat), .Y(G3280GAT_1144_gat) );
AND2XL U_g1114 (.A(G3157GAT_1101_ngat), .B(G3221GAT_1124_ngat), .Y(G3276GAT_1145_gat) );
AND2XL U_g1115 (.A(G3152GAT_1103_ngat), .B(G3218GAT_1125_ngat), .Y(G3272GAT_1146_gat) );
AND2XL U_g1116 (.A(G3147GAT_1105_ngat), .B(G3215GAT_1126_ngat), .Y(G3268GAT_1147_gat) );
AND2XL U_g1117 (.A(G3142GAT_1107_ngat), .B(G3212GAT_1127_ngat), .Y(G3264GAT_1148_gat) );
AND2XL U_g1118 (.A(G3322GAT_1130_ngat), .B(G3321GAT_1129_ngat), .Y(G3362GAT_1149_gat) );
AND2XL U_g1119 (.A(G3317GAT_1131_ngat), .B(G3257GAT_1110_ngat), .Y(G3360GAT_1150_gat) );
AND2XL U_g1120 (.A(G3254GAT_1111_ngat), .B(G3317GAT_1131_ngat), .Y(G3361GAT_1151_gat) );
AND2XL U_g1121 (.A(G3311GAT_1133_ngat), .B(G3314GAT_1132_ngat), .Y(G3356GAT_1152_gat) );
AND2XL U_g1122 (.A(G3310GAT_1137_ngat), .B(G3309GAT_1134_ngat), .Y(G3353GAT_1153_gat) );
AND2XL U_g1123 (.A(G3305GAT_1138_ngat), .B(G3127GAT_1054_ngat), .Y(G3350GAT_1154_gat) );
AND2XL U_g1124 (.A(G3305GAT_1138_ngat), .B(G3245GAT_1113_ngat), .Y(G3348GAT_1155_gat) );
AND2XL U_g1125 (.A(G3301GAT_1139_ngat), .B(G3300GAT_1136_ngat), .Y(G3341GAT_1156_gat) );
AND2XL U_g1126 (.A(G3296GAT_1140_ngat), .B(G3236GAT_1117_ngat), .Y(G3339GAT_1157_gat) );
AND2XL U_g1127 (.A(G3292GAT_1141_ngat), .B(G3233GAT_1118_ngat), .Y(G3337GAT_1158_gat) );
AND2XL U_g1128 (.A(G3288GAT_1142_ngat), .B(G3230GAT_1120_ngat), .Y(G3335GAT_1159_gat) );
AND2XL U_g1129 (.A(G3284GAT_1143_ngat), .B(G3227GAT_1122_ngat), .Y(G3333GAT_1160_gat) );
AND2XL U_g1130 (.A(G1092GAT_104_ngat), .B(G3305GAT_1138_ngat), .Y(G3349GAT_1161_gat) );
AND2XL U_g1131 (.A(G3280GAT_1144_ngat), .B(G3224GAT_1123_ngat), .Y(G3331GAT_1162_gat) );
AND2XL U_g1132 (.A(G1044GAT_120_ngat), .B(G3302GAT_1135_ngat), .Y(G3344GAT_1163_gat) );
AND2XL U_g1133 (.A(G3276GAT_1145_ngat), .B(G3221GAT_1124_ngat), .Y(G3329GAT_1164_gat) );
AND2XL U_g1134 (.A(G3182GAT_1087_ngat), .B(G3296GAT_1140_ngat), .Y(G3340GAT_1165_gat) );
AND2XL U_g1135 (.A(G3272GAT_1146_ngat), .B(G3218GAT_1125_ngat), .Y(G3327GAT_1166_gat) );
AND2XL U_g1136 (.A(G3177GAT_1090_ngat), .B(G3292GAT_1141_ngat), .Y(G3338GAT_1167_gat) );
AND2XL U_g1137 (.A(G3268GAT_1147_ngat), .B(G3215GAT_1126_ngat), .Y(G3325GAT_1168_gat) );
AND2XL U_g1138 (.A(G3172GAT_1093_ngat), .B(G3288GAT_1142_ngat), .Y(G3336GAT_1169_gat) );
AND2XL U_g1139 (.A(G3264GAT_1148_ngat), .B(G3212GAT_1127_ngat), .Y(G3323GAT_1170_gat) );
AND2XL U_g1140 (.A(G3167GAT_1096_ngat), .B(G3284GAT_1143_ngat), .Y(G3334GAT_1171_gat) );
AND2XL U_g1141 (.A(G3162GAT_1099_ngat), .B(G3280GAT_1144_ngat), .Y(G3332GAT_1172_gat) );
AND2XL U_g1142 (.A(G3157GAT_1101_ngat), .B(G3276GAT_1145_ngat), .Y(G3330GAT_1173_gat) );
AND2XL U_g1143 (.A(G3152GAT_1103_ngat), .B(G3272GAT_1146_ngat), .Y(G3328GAT_1174_gat) );
AND2XL U_g1144 (.A(G3147GAT_1105_ngat), .B(G3268GAT_1147_ngat), .Y(G3326GAT_1175_gat) );
AND2XL U_g1145 (.A(G3142GAT_1107_ngat), .B(G3264GAT_1148_ngat), .Y(G3324GAT_1176_gat) );
AND2XL U_g1146 (.A(G3361GAT_1151_ngat), .B(G3360GAT_1150_ngat), .Y(G3410GAT_1177_gat) );
AND2XL U_g1147 (.A(G3356GAT_1152_ngat), .B(G3314GAT_1132_ngat), .Y(G3408GAT_1178_gat) );
AND2XL U_g1148 (.A(G3311GAT_1133_ngat), .B(G3356GAT_1152_ngat), .Y(G3409GAT_1179_gat) );
AND2XL U_g1149 (.A(G3350GAT_1154_ngat), .B(G3353GAT_1153_ngat), .Y(G3404GAT_1180_gat) );
AND2XL U_g1150 (.A(G3349GAT_1161_ngat), .B(G3348GAT_1155_ngat), .Y(G3401GAT_1181_gat) );
AND2XL U_g1151 (.A(G3344GAT_1163_ngat), .B(G3193GAT_1075_ngat), .Y(G3398GAT_1182_gat) );
AND2XL U_g1152 (.A(G3344GAT_1163_ngat), .B(G3302GAT_1135_ngat), .Y(G3396GAT_1183_gat) );
AND2XL U_g1153 (.A(G3340GAT_1165_ngat), .B(G3339GAT_1157_ngat), .Y(G3389GAT_1184_gat) );
AND2XL U_g1154 (.A(G1239GAT_55_ngat), .B(G3362GAT_1149_ngat), .Y(G3413GAT_1185_gat) );
AND2XL U_g1155 (.A(G3338GAT_1167_ngat), .B(G3337GAT_1158_ngat), .Y(G3386GAT_1186_gat) );
AND2XL U_g1156 (.A(G3336GAT_1169_ngat), .B(G3335GAT_1159_ngat), .Y(G3383GAT_1187_gat) );
AND2XL U_g1157 (.A(G3334GAT_1171_ngat), .B(G3333GAT_1160_ngat), .Y(G3380GAT_1188_gat) );
AND2XL U_g1158 (.A(G3332GAT_1172_ngat), .B(G3331GAT_1162_ngat), .Y(G3377GAT_1189_gat) );
AND2XL U_g1159 (.A(G1044GAT_120_ngat), .B(G3344GAT_1163_ngat), .Y(G3397GAT_1190_gat) );
AND2XL U_g1160 (.A(G3330GAT_1173_ngat), .B(G3329GAT_1164_ngat), .Y(G3374GAT_1191_gat) );
AND2XL U_g1161 (.A(G996GAT_136_ngat), .B(G3341GAT_1156_ngat), .Y(G3392GAT_1192_gat) );
AND2XL U_g1162 (.A(G3328GAT_1174_ngat), .B(G3327GAT_1166_ngat), .Y(G3371GAT_1193_gat) );
AND2XL U_g1163 (.A(G3326GAT_1175_ngat), .B(G3325GAT_1168_ngat), .Y(G3368GAT_1194_gat) );
AND2XL U_g1164 (.A(G3324GAT_1176_ngat), .B(G3323GAT_1170_ngat), .Y(G3365GAT_1195_gat) );
AND2XL U_g1165 (.A(G3413GAT_1185_ngat), .B(G3260GAT_1109_ngat), .Y(G3476GAT_1196_gat) );
AND2XL U_g1166 (.A(G3413GAT_1185_ngat), .B(G3362GAT_1149_ngat), .Y(G3474GAT_1197_gat) );
AND2XL U_g1167 (.A(G3409GAT_1179_ngat), .B(G3408GAT_1178_ngat), .Y(G3467GAT_1198_gat) );
AND2XL U_g1168 (.A(G3404GAT_1180_ngat), .B(G3353GAT_1153_ngat), .Y(G3465GAT_1199_gat) );
AND2XL U_g1169 (.A(G3350GAT_1154_ngat), .B(G3404GAT_1180_ngat), .Y(G3466GAT_1200_gat) );
AND2XL U_g1170 (.A(G3398GAT_1182_ngat), .B(G3401GAT_1181_ngat), .Y(G3461GAT_1201_gat) );
AND2XL U_g1171 (.A(G3397GAT_1190_ngat), .B(G3396GAT_1183_ngat), .Y(G3458GAT_1202_gat) );
AND2XL U_g1172 (.A(G3392GAT_1192_ngat), .B(G3239GAT_1116_ngat), .Y(G3455GAT_1203_gat) );
AND2XL U_g1173 (.A(G3392GAT_1192_ngat), .B(G3341GAT_1156_ngat), .Y(G3453GAT_1204_gat) );
AND2XL U_g1174 (.A(G1239GAT_55_ngat), .B(G3413GAT_1185_ngat), .Y(G3475GAT_1205_gat) );
AND2XL U_g1175 (.A(G1191GAT_71_ngat), .B(G3410GAT_1177_ngat), .Y(G3470GAT_1206_gat) );
AND2XL U_g1176 (.A(G996GAT_136_ngat), .B(G3392GAT_1192_ngat), .Y(G3454GAT_1207_gat) );
AND2XL U_g1177 (.A(G948GAT_152_ngat), .B(G3389GAT_1184_ngat), .Y(G3449GAT_1208_gat) );
AND2XL U_g1178 (.A(G900GAT_168_ngat), .B(G3386GAT_1186_ngat), .Y(G3445GAT_1209_gat) );
AND2XL U_g1179 (.A(G852GAT_184_ngat), .B(G3383GAT_1187_ngat), .Y(G3441GAT_1210_gat) );
AND2XL U_g1180 (.A(G804GAT_200_ngat), .B(G3380GAT_1188_ngat), .Y(G3437GAT_1211_gat) );
AND2XL U_g1181 (.A(G756GAT_216_ngat), .B(G3377GAT_1189_ngat), .Y(G3433GAT_1212_gat) );
AND2XL U_g1182 (.A(G708GAT_232_ngat), .B(G3374GAT_1191_ngat), .Y(G3429GAT_1213_gat) );
AND2XL U_g1183 (.A(G660GAT_248_ngat), .B(G3371GAT_1193_ngat), .Y(G3425GAT_1214_gat) );
AND2XL U_g1184 (.A(G612GAT_264_ngat), .B(G3368GAT_1194_ngat), .Y(G3421GAT_1215_gat) );
AND2XL U_g1185 (.A(G564GAT_280_ngat), .B(G3365GAT_1195_ngat), .Y(G3417GAT_1216_gat) );
AND2XL U_g1186 (.A(G3476GAT_1196_ngat), .B(G1287GAT_39_ngat), .Y(G3548GAT_1217_gat) );
AND2XL U_g1187 (.A(G3475GAT_1205_ngat), .B(G3474GAT_1197_ngat), .Y(G3545GAT_1218_gat) );
AND2XL U_g1188 (.A(G3470GAT_1206_ngat), .B(G3317GAT_1131_ngat), .Y(G3542GAT_1219_gat) );
AND2XL U_g1189 (.A(G3470GAT_1206_ngat), .B(G3410GAT_1177_ngat), .Y(G3540GAT_1220_gat) );
AND2XL U_g1190 (.A(G3466GAT_1200_ngat), .B(G3465GAT_1199_ngat), .Y(G3533GAT_1221_gat) );
AND2XL U_g1191 (.A(G3461GAT_1201_ngat), .B(G3401GAT_1181_ngat), .Y(G3531GAT_1222_gat) );
AND2XL U_g1192 (.A(G3398GAT_1182_ngat), .B(G3461GAT_1201_ngat), .Y(G3532GAT_1223_gat) );
AND2XL U_g1193 (.A(G3455GAT_1203_ngat), .B(G3458GAT_1202_ngat), .Y(G3527GAT_1224_gat) );
AND2XL U_g1194 (.A(G3454GAT_1207_ngat), .B(G3453GAT_1204_ngat), .Y(G3524GAT_1225_gat) );
AND2XL U_g1195 (.A(G3449GAT_1208_ngat), .B(G3389GAT_1184_ngat), .Y(G3519GAT_1226_gat) );
AND2XL U_g1196 (.A(G3445GAT_1209_ngat), .B(G3386GAT_1186_ngat), .Y(G3514GAT_1227_gat) );
AND2XL U_g1197 (.A(G1191GAT_71_ngat), .B(G3470GAT_1206_ngat), .Y(G3541GAT_1228_gat) );
AND2XL U_g1198 (.A(G3441GAT_1210_ngat), .B(G3383GAT_1187_ngat), .Y(G3509GAT_1229_gat) );
AND2XL U_g1199 (.A(G1143GAT_87_ngat), .B(G3467GAT_1198_ngat), .Y(G3536GAT_1230_gat) );
AND2XL U_g1200 (.A(G3437GAT_1211_ngat), .B(G3380GAT_1188_ngat), .Y(G3504GAT_1231_gat) );
AND2XL U_g1201 (.A(G3433GAT_1212_ngat), .B(G3377GAT_1189_ngat), .Y(G3499GAT_1232_gat) );
AND2XL U_g1202 (.A(G3429GAT_1213_ngat), .B(G3374GAT_1191_ngat), .Y(G3494GAT_1233_gat) );
AND2XL U_g1203 (.A(G3449GAT_1208_ngat), .B(G3296GAT_1140_ngat), .Y(G3521GAT_1234_gat) );
AND2XL U_g1204 (.A(G3425GAT_1214_ngat), .B(G3371GAT_1193_ngat), .Y(G3489GAT_1235_gat) );
AND2XL U_g1205 (.A(G948GAT_152_ngat), .B(G3449GAT_1208_ngat), .Y(G3520GAT_1236_gat) );
AND2XL U_g1206 (.A(G3445GAT_1209_ngat), .B(G3292GAT_1141_ngat), .Y(G3516GAT_1237_gat) );
AND2XL U_g1207 (.A(G3421GAT_1215_ngat), .B(G3368GAT_1194_ngat), .Y(G3484GAT_1238_gat) );
AND2XL U_g1208 (.A(G900GAT_168_ngat), .B(G3445GAT_1209_ngat), .Y(G3515GAT_1239_gat) );
AND2XL U_g1209 (.A(G3441GAT_1210_ngat), .B(G3288GAT_1142_ngat), .Y(G3511GAT_1240_gat) );
AND2XL U_g1210 (.A(G3417GAT_1216_ngat), .B(G3365GAT_1195_ngat), .Y(G3479GAT_1241_gat) );
AND2XL U_g1211 (.A(G852GAT_184_ngat), .B(G3441GAT_1210_ngat), .Y(G3510GAT_1242_gat) );
AND2XL U_g1212 (.A(G3437GAT_1211_ngat), .B(G3284GAT_1143_ngat), .Y(G3506GAT_1243_gat) );
AND2XL U_g1213 (.A(G804GAT_200_ngat), .B(G3437GAT_1211_ngat), .Y(G3505GAT_1244_gat) );
AND2XL U_g1214 (.A(G3433GAT_1212_ngat), .B(G3280GAT_1144_ngat), .Y(G3501GAT_1245_gat) );
AND2XL U_g1215 (.A(G756GAT_216_ngat), .B(G3433GAT_1212_ngat), .Y(G3500GAT_1246_gat) );
AND2XL U_g1216 (.A(G3429GAT_1213_ngat), .B(G3276GAT_1145_ngat), .Y(G3496GAT_1247_gat) );
AND2XL U_g1217 (.A(G708GAT_232_ngat), .B(G3429GAT_1213_ngat), .Y(G3495GAT_1248_gat) );
AND2XL U_g1218 (.A(G3425GAT_1214_ngat), .B(G3272GAT_1146_ngat), .Y(G3491GAT_1249_gat) );
AND2XL U_g1219 (.A(G660GAT_248_ngat), .B(G3425GAT_1214_ngat), .Y(G3490GAT_1250_gat) );
AND2XL U_g1220 (.A(G3421GAT_1215_ngat), .B(G3268GAT_1147_ngat), .Y(G3486GAT_1251_gat) );
AND2XL U_g1221 (.A(G612GAT_264_ngat), .B(G3421GAT_1215_ngat), .Y(G3485GAT_1252_gat) );
AND2XL U_g1222 (.A(G3417GAT_1216_ngat), .B(G3264GAT_1148_ngat), .Y(G3481GAT_1253_gat) );
AND2XL U_g1223 (.A(G564GAT_280_ngat), .B(G3417GAT_1216_ngat), .Y(G3480GAT_1254_gat) );
AND2XL U_g1224 (.A(G3548GAT_1217_ngat), .B(G1287GAT_39_ngat), .Y(G3602GAT_1255_gat) );
AND2XL U_g1225 (.A(G3476GAT_1196_ngat), .B(G3548GAT_1217_ngat), .Y(G3603GAT_1256_gat) );
AND2XL U_g1226 (.A(G3542GAT_1219_ngat), .B(G3545GAT_1218_ngat), .Y(G3598GAT_1257_gat) );
AND2XL U_g1227 (.A(G3541GAT_1228_ngat), .B(G3540GAT_1220_ngat), .Y(G3595GAT_1258_gat) );
AND2XL U_g1228 (.A(G3536GAT_1230_ngat), .B(G3356GAT_1152_ngat), .Y(G3592GAT_1259_gat) );
AND2XL U_g1229 (.A(G3536GAT_1230_ngat), .B(G3467GAT_1198_ngat), .Y(G3590GAT_1260_gat) );
AND2XL U_g1230 (.A(G3532GAT_1223_ngat), .B(G3531GAT_1222_ngat), .Y(G3583GAT_1261_gat) );
AND2XL U_g1231 (.A(G3527GAT_1224_ngat), .B(G3458GAT_1202_ngat), .Y(G3581GAT_1262_gat) );
AND2XL U_g1232 (.A(G3455GAT_1203_ngat), .B(G3527GAT_1224_ngat), .Y(G3582GAT_1263_gat) );
AND2XL U_g1233 (.A(G3521GAT_1234_ngat), .B(G3524GAT_1225_ngat), .Y(G3577GAT_1264_gat) );
AND2XL U_g1234 (.A(G3520GAT_1236_ngat), .B(G3519GAT_1226_ngat), .Y(G3574GAT_1265_gat) );
AND2XL U_g1235 (.A(G3515GAT_1239_ngat), .B(G3514GAT_1227_ngat), .Y(G3571GAT_1266_gat) );
AND2XL U_g1236 (.A(G3510GAT_1242_ngat), .B(G3509GAT_1229_ngat), .Y(G3568GAT_1267_gat) );
AND2XL U_g1237 (.A(G1143GAT_87_ngat), .B(G3536GAT_1230_ngat), .Y(G3591GAT_1268_gat) );
AND2XL U_g1238 (.A(G3505GAT_1244_ngat), .B(G3504GAT_1231_ngat), .Y(G3565GAT_1269_gat) );
AND2XL U_g1239 (.A(G1095GAT_103_ngat), .B(G3533GAT_1221_ngat), .Y(G3586GAT_1270_gat) );
AND2XL U_g1240 (.A(G3500GAT_1246_ngat), .B(G3499GAT_1232_ngat), .Y(G3562GAT_1271_gat) );
AND2XL U_g1241 (.A(G3495GAT_1248_ngat), .B(G3494GAT_1233_ngat), .Y(G3559GAT_1272_gat) );
AND2XL U_g1242 (.A(G3490GAT_1250_ngat), .B(G3489GAT_1235_ngat), .Y(G3556GAT_1273_gat) );
AND2XL U_g1243 (.A(G3485GAT_1252_ngat), .B(G3484GAT_1238_ngat), .Y(G3553GAT_1274_gat) );
AND2XL U_g1244 (.A(G3480GAT_1254_ngat), .B(G3479GAT_1241_ngat), .Y(G3552GAT_1275_gat) );
AND2XL U_g1245 (.A(G3603GAT_1256_ngat), .B(G3602GAT_1255_ngat), .Y(G3659GAT_1276_gat) );
AND2XL U_g1246 (.A(G3598GAT_1257_ngat), .B(G3545GAT_1218_ngat), .Y(G3657GAT_1277_gat) );
AND2XL U_g1247 (.A(G3542GAT_1219_ngat), .B(G3598GAT_1257_ngat), .Y(G3658GAT_1278_gat) );
AND2XL U_g1248 (.A(G3592GAT_1259_ngat), .B(G3595GAT_1258_ngat), .Y(G3653GAT_1279_gat) );
AND2XL U_g1249 (.A(G3591GAT_1268_ngat), .B(G3590GAT_1260_ngat), .Y(G3650GAT_1280_gat) );
AND2XL U_g1250 (.A(G3586GAT_1270_ngat), .B(G3404GAT_1180_ngat), .Y(G3647GAT_1281_gat) );
AND2XL U_g1251 (.A(G3586GAT_1270_ngat), .B(G3533GAT_1221_ngat), .Y(G3645GAT_1282_gat) );
AND2XL U_g1252 (.A(G3582GAT_1263_ngat), .B(G3581GAT_1262_ngat), .Y(G3638GAT_1283_gat) );
AND2XL U_g1253 (.A(G3577GAT_1264_ngat), .B(G3524GAT_1225_ngat), .Y(G3636GAT_1284_gat) );
AND2XL U_g1254 (.A(G1095GAT_103_ngat), .B(G3586GAT_1270_ngat), .Y(G3646GAT_1285_gat) );
AND2XL U_g1255 (.A(G1047GAT_119_ngat), .B(G3583GAT_1261_ngat), .Y(G3641GAT_1286_gat) );
AND2XL U_g1256 (.A(G3521GAT_1234_ngat), .B(G3577GAT_1264_ngat), .Y(G3637GAT_1287_gat) );
AND2XL U_g1257 (.A(G3516GAT_1237_ngat), .B(G3574GAT_1265_ngat), .Y(G3632GAT_1288_gat) );
AND2XL U_g1258 (.A(G3511GAT_1240_ngat), .B(G3571GAT_1266_ngat), .Y(G3628GAT_1289_gat) );
AND2XL U_g1259 (.A(G3506GAT_1243_ngat), .B(G3568GAT_1267_ngat), .Y(G3624GAT_1290_gat) );
AND2XL U_g1260 (.A(G3501GAT_1245_ngat), .B(G3565GAT_1269_ngat), .Y(G3620GAT_1291_gat) );
AND2XL U_g1261 (.A(G3496GAT_1247_ngat), .B(G3562GAT_1271_ngat), .Y(G3616GAT_1292_gat) );
AND2XL U_g1262 (.A(G3491GAT_1249_ngat), .B(G3559GAT_1272_ngat), .Y(G3612GAT_1293_gat) );
AND2XL U_g1263 (.A(G3486GAT_1251_ngat), .B(G3556GAT_1273_ngat), .Y(G3608GAT_1294_gat) );
AND2XL U_g1264 (.A(G3481GAT_1253_ngat), .B(G3553GAT_1274_ngat), .Y(G3604GAT_1295_gat) );
AND2XL U_g1265 (.A(G3658GAT_1278_ngat), .B(G3657GAT_1277_ngat), .Y(G3699GAT_1296_gat) );
AND2XL U_g1266 (.A(G3653GAT_1279_ngat), .B(G3595GAT_1258_ngat), .Y(G3697GAT_1297_gat) );
AND2XL U_g1267 (.A(G3592GAT_1259_ngat), .B(G3653GAT_1279_ngat), .Y(G3698GAT_1298_gat) );
AND2XL U_g1268 (.A(G3647GAT_1281_ngat), .B(G3650GAT_1280_ngat), .Y(G3693GAT_1299_gat) );
AND2XL U_g1269 (.A(G3646GAT_1285_ngat), .B(G3645GAT_1282_ngat), .Y(G3690GAT_1300_gat) );
AND2XL U_g1270 (.A(G3641GAT_1286_ngat), .B(G3461GAT_1201_ngat), .Y(G3687GAT_1301_gat) );
AND2XL U_g1271 (.A(G3641GAT_1286_ngat), .B(G3583GAT_1261_ngat), .Y(G3685GAT_1302_gat) );
AND2XL U_g1272 (.A(G3637GAT_1287_ngat), .B(G3636GAT_1284_ngat), .Y(G3678GAT_1303_gat) );
AND2XL U_g1273 (.A(G3632GAT_1288_ngat), .B(G3574GAT_1265_ngat), .Y(G3676GAT_1304_gat) );
AND2XL U_g1274 (.A(G1242GAT_54_ngat), .B(G3659GAT_1276_ngat), .Y(G3702GAT_1305_gat) );
AND2XL U_g1275 (.A(G3628GAT_1289_ngat), .B(G3571GAT_1266_ngat), .Y(G3674GAT_1306_gat) );
AND2XL U_g1276 (.A(G3624GAT_1290_ngat), .B(G3568GAT_1267_ngat), .Y(G3672GAT_1307_gat) );
AND2XL U_g1277 (.A(G3620GAT_1291_ngat), .B(G3565GAT_1269_ngat), .Y(G3670GAT_1308_gat) );
AND2XL U_g1278 (.A(G3616GAT_1292_ngat), .B(G3562GAT_1271_ngat), .Y(G3668GAT_1309_gat) );
AND2XL U_g1279 (.A(G1047GAT_119_ngat), .B(G3641GAT_1286_ngat), .Y(G3686GAT_1310_gat) );
AND2XL U_g1280 (.A(G3612GAT_1293_ngat), .B(G3559GAT_1272_ngat), .Y(G3666GAT_1311_gat) );
AND2XL U_g1281 (.A(G999GAT_135_ngat), .B(G3638GAT_1283_ngat), .Y(G3681GAT_1312_gat) );
AND2XL U_g1282 (.A(G3608GAT_1294_ngat), .B(G3556GAT_1273_ngat), .Y(G3664GAT_1313_gat) );
AND2XL U_g1283 (.A(G3516GAT_1237_ngat), .B(G3632GAT_1288_ngat), .Y(G3677GAT_1314_gat) );
AND2XL U_g1284 (.A(G3604GAT_1295_ngat), .B(G3553GAT_1274_ngat), .Y(G3662GAT_1315_gat) );
AND2XL U_g1285 (.A(G3511GAT_1240_ngat), .B(G3628GAT_1289_ngat), .Y(G3675GAT_1316_gat) );
AND2XL U_g1286 (.A(G3506GAT_1243_ngat), .B(G3624GAT_1290_ngat), .Y(G3673GAT_1317_gat) );
AND2XL U_g1287 (.A(G3501GAT_1245_ngat), .B(G3620GAT_1291_ngat), .Y(G3671GAT_1318_gat) );
AND2XL U_g1288 (.A(G3496GAT_1247_ngat), .B(G3616GAT_1292_ngat), .Y(G3669GAT_1319_gat) );
AND2XL U_g1289 (.A(G3491GAT_1249_ngat), .B(G3612GAT_1293_ngat), .Y(G3667GAT_1320_gat) );
AND2XL U_g1290 (.A(G3486GAT_1251_ngat), .B(G3608GAT_1294_ngat), .Y(G3665GAT_1321_gat) );
AND2XL U_g1291 (.A(G3481GAT_1253_ngat), .B(G3604GAT_1295_ngat), .Y(G3663GAT_1322_gat) );
AND2XL U_g1292 (.A(G3702GAT_1305_ngat), .B(G3548GAT_1217_ngat), .Y(G3757GAT_1323_gat) );
AND2XL U_g1293 (.A(G3702GAT_1305_ngat), .B(G3659GAT_1276_ngat), .Y(G3755GAT_1324_gat) );
AND2XL U_g1294 (.A(G3698GAT_1298_ngat), .B(G3697GAT_1297_ngat), .Y(G3748GAT_1325_gat) );
AND2XL U_g1295 (.A(G3693GAT_1299_ngat), .B(G3650GAT_1280_ngat), .Y(G3746GAT_1326_gat) );
AND2XL U_g1296 (.A(G3647GAT_1281_ngat), .B(G3693GAT_1299_ngat), .Y(G3747GAT_1327_gat) );
AND2XL U_g1297 (.A(G3687GAT_1301_ngat), .B(G3690GAT_1300_ngat), .Y(G3742GAT_1328_gat) );
AND2XL U_g1298 (.A(G3686GAT_1310_ngat), .B(G3685GAT_1302_ngat), .Y(G3739GAT_1329_gat) );
AND2XL U_g1299 (.A(G3681GAT_1312_ngat), .B(G3527GAT_1224_ngat), .Y(G3736GAT_1330_gat) );
AND2XL U_g1300 (.A(G3681GAT_1312_ngat), .B(G3638GAT_1283_ngat), .Y(G3734GAT_1331_gat) );
AND2XL U_g1301 (.A(G3677GAT_1314_ngat), .B(G3676GAT_1304_ngat), .Y(G3727GAT_1332_gat) );
AND2XL U_g1302 (.A(G1242GAT_54_ngat), .B(G3702GAT_1305_ngat), .Y(G3756GAT_1333_gat) );
AND2XL U_g1303 (.A(G3675GAT_1316_ngat), .B(G3674GAT_1306_ngat), .Y(G3724GAT_1334_gat) );
AND2XL U_g1304 (.A(G1194GAT_70_ngat), .B(G3699GAT_1296_ngat), .Y(G3751GAT_1335_gat) );
AND2XL U_g1305 (.A(G3673GAT_1317_ngat), .B(G3672GAT_1307_ngat), .Y(G3721GAT_1336_gat) );
AND2XL U_g1306 (.A(G3671GAT_1318_ngat), .B(G3670GAT_1308_ngat), .Y(G3718GAT_1337_gat) );
AND2XL U_g1307 (.A(G3669GAT_1319_ngat), .B(G3668GAT_1309_ngat), .Y(G3715GAT_1338_gat) );
AND2XL U_g1308 (.A(G3667GAT_1320_ngat), .B(G3666GAT_1311_ngat), .Y(G3712GAT_1339_gat) );
AND2XL U_g1309 (.A(G999GAT_135_ngat), .B(G3681GAT_1312_ngat), .Y(G3735GAT_1340_gat) );
AND2XL U_g1310 (.A(G3665GAT_1321_ngat), .B(G3664GAT_1313_ngat), .Y(G3709GAT_1341_gat) );
AND2XL U_g1311 (.A(G951GAT_151_ngat), .B(G3678GAT_1303_ngat), .Y(G3730GAT_1342_gat) );
AND2XL U_g1312 (.A(G3663GAT_1322_ngat), .B(G3662GAT_1315_ngat), .Y(G3706GAT_1343_gat) );
AND2XL U_g1313 (.A(G3757GAT_1323_ngat), .B(G1290GAT_38_ngat), .Y(G3821GAT_1344_gat) );
AND2XL U_g1314 (.A(G3756GAT_1333_ngat), .B(G3755GAT_1324_ngat), .Y(G3818GAT_1345_gat) );
AND2XL U_g1315 (.A(G3751GAT_1335_ngat), .B(G3598GAT_1257_ngat), .Y(G3815GAT_1346_gat) );
AND2XL U_g1316 (.A(G3751GAT_1335_ngat), .B(G3699GAT_1296_ngat), .Y(G3813GAT_1347_gat) );
AND2XL U_g1317 (.A(G3747GAT_1327_ngat), .B(G3746GAT_1326_ngat), .Y(G3806GAT_1348_gat) );
AND2XL U_g1318 (.A(G3742GAT_1328_ngat), .B(G3690GAT_1300_ngat), .Y(G3804GAT_1349_gat) );
AND2XL U_g1319 (.A(G3687GAT_1301_ngat), .B(G3742GAT_1328_ngat), .Y(G3805GAT_1350_gat) );
AND2XL U_g1320 (.A(G3736GAT_1330_ngat), .B(G3739GAT_1329_ngat), .Y(G3800GAT_1351_gat) );
AND2XL U_g1321 (.A(G3735GAT_1340_ngat), .B(G3734GAT_1331_ngat), .Y(G3797GAT_1352_gat) );
AND2XL U_g1322 (.A(G3730GAT_1342_ngat), .B(G3577GAT_1264_ngat), .Y(G3794GAT_1353_gat) );
AND2XL U_g1323 (.A(G3730GAT_1342_ngat), .B(G3678GAT_1303_ngat), .Y(G3792GAT_1354_gat) );
AND2XL U_g1324 (.A(G1194GAT_70_ngat), .B(G3751GAT_1335_ngat), .Y(G3814GAT_1355_gat) );
AND2XL U_g1325 (.A(G1146GAT_86_ngat), .B(G3748GAT_1325_ngat), .Y(G3809GAT_1356_gat) );
AND2XL U_g1326 (.A(G951GAT_151_ngat), .B(G3730GAT_1342_ngat), .Y(G3793GAT_1357_gat) );
AND2XL U_g1327 (.A(G903GAT_167_ngat), .B(G3727GAT_1332_ngat), .Y(G3788GAT_1358_gat) );
AND2XL U_g1328 (.A(G855GAT_183_ngat), .B(G3724GAT_1334_ngat), .Y(G3784GAT_1359_gat) );
AND2XL U_g1329 (.A(G807GAT_199_ngat), .B(G3721GAT_1336_ngat), .Y(G3780GAT_1360_gat) );
AND2XL U_g1330 (.A(G759GAT_215_ngat), .B(G3718GAT_1337_ngat), .Y(G3776GAT_1361_gat) );
AND2XL U_g1331 (.A(G711GAT_231_ngat), .B(G3715GAT_1338_ngat), .Y(G3772GAT_1362_gat) );
AND2XL U_g1332 (.A(G663GAT_247_ngat), .B(G3712GAT_1339_ngat), .Y(G3768GAT_1363_gat) );
AND2XL U_g1333 (.A(G615GAT_263_ngat), .B(G3709GAT_1341_ngat), .Y(G3764GAT_1364_gat) );
AND2XL U_g1334 (.A(G567GAT_279_ngat), .B(G3706GAT_1343_ngat), .Y(G3760GAT_1365_gat) );
AND2XL U_g1335 (.A(G3821GAT_1344_ngat), .B(G1290GAT_38_ngat), .Y(G3893GAT_1366_gat) );
AND2XL U_g1336 (.A(G3757GAT_1323_ngat), .B(G3821GAT_1344_ngat), .Y(G3894GAT_1367_gat) );
AND2XL U_g1337 (.A(G3815GAT_1346_ngat), .B(G3818GAT_1345_ngat), .Y(G3889GAT_1368_gat) );
AND2XL U_g1338 (.A(G3814GAT_1355_ngat), .B(G3813GAT_1347_ngat), .Y(G3886GAT_1369_gat) );
AND2XL U_g1339 (.A(G3809GAT_1356_ngat), .B(G3653GAT_1279_ngat), .Y(G3883GAT_1370_gat) );
AND2XL U_g1340 (.A(G3809GAT_1356_ngat), .B(G3748GAT_1325_ngat), .Y(G3881GAT_1371_gat) );
AND2XL U_g1341 (.A(G3805GAT_1350_ngat), .B(G3804GAT_1349_ngat), .Y(G3874GAT_1372_gat) );
AND2XL U_g1342 (.A(G3800GAT_1351_ngat), .B(G3739GAT_1329_ngat), .Y(G3872GAT_1373_gat) );
AND2XL U_g1343 (.A(G3736GAT_1330_ngat), .B(G3800GAT_1351_ngat), .Y(G3873GAT_1374_gat) );
AND2XL U_g1344 (.A(G3794GAT_1353_ngat), .B(G3797GAT_1352_ngat), .Y(G3868GAT_1375_gat) );
AND2XL U_g1345 (.A(G3793GAT_1357_ngat), .B(G3792GAT_1354_ngat), .Y(G3865GAT_1376_gat) );
AND2XL U_g1346 (.A(G3788GAT_1358_ngat), .B(G3727GAT_1332_ngat), .Y(G3860GAT_1377_gat) );
AND2XL U_g1347 (.A(G3784GAT_1359_ngat), .B(G3724GAT_1334_ngat), .Y(G3855GAT_1378_gat) );
AND2XL U_g1348 (.A(G3780GAT_1360_ngat), .B(G3721GAT_1336_ngat), .Y(G3850GAT_1379_gat) );
AND2XL U_g1349 (.A(G1146GAT_86_ngat), .B(G3809GAT_1356_ngat), .Y(G3882GAT_1380_gat) );
AND2XL U_g1350 (.A(G3776GAT_1361_ngat), .B(G3718GAT_1337_ngat), .Y(G3845GAT_1381_gat) );
AND2XL U_g1351 (.A(G1098GAT_102_ngat), .B(G3806GAT_1348_ngat), .Y(G3877GAT_1382_gat) );
AND2XL U_g1352 (.A(G3772GAT_1362_ngat), .B(G3715GAT_1338_ngat), .Y(G3840GAT_1383_gat) );
AND2XL U_g1353 (.A(G3768GAT_1363_ngat), .B(G3712GAT_1339_ngat), .Y(G3835GAT_1384_gat) );
AND2XL U_g1354 (.A(G3764GAT_1364_ngat), .B(G3709GAT_1341_ngat), .Y(G3830GAT_1385_gat) );
AND2XL U_g1355 (.A(G3788GAT_1358_ngat), .B(G3632GAT_1288_ngat), .Y(G3862GAT_1386_gat) );
AND2XL U_g1356 (.A(G3760GAT_1365_ngat), .B(G3706GAT_1343_ngat), .Y(G3825GAT_1387_gat) );
AND2XL U_g1357 (.A(G903GAT_167_ngat), .B(G3788GAT_1358_ngat), .Y(G3861GAT_1388_gat) );
AND2XL U_g1358 (.A(G3784GAT_1359_ngat), .B(G3628GAT_1289_ngat), .Y(G3857GAT_1389_gat) );
AND2XL U_g1359 (.A(G855GAT_183_ngat), .B(G3784GAT_1359_ngat), .Y(G3856GAT_1390_gat) );
AND2XL U_g1360 (.A(G3780GAT_1360_ngat), .B(G3624GAT_1290_ngat), .Y(G3852GAT_1391_gat) );
AND2XL U_g1361 (.A(G807GAT_199_ngat), .B(G3780GAT_1360_ngat), .Y(G3851GAT_1392_gat) );
AND2XL U_g1362 (.A(G3776GAT_1361_ngat), .B(G3620GAT_1291_ngat), .Y(G3847GAT_1393_gat) );
AND2XL U_g1363 (.A(G759GAT_215_ngat), .B(G3776GAT_1361_ngat), .Y(G3846GAT_1394_gat) );
AND2XL U_g1364 (.A(G3772GAT_1362_ngat), .B(G3616GAT_1292_ngat), .Y(G3842GAT_1395_gat) );
AND2XL U_g1365 (.A(G711GAT_231_ngat), .B(G3772GAT_1362_ngat), .Y(G3841GAT_1396_gat) );
AND2XL U_g1366 (.A(G3768GAT_1363_ngat), .B(G3612GAT_1293_ngat), .Y(G3837GAT_1397_gat) );
AND2XL U_g1367 (.A(G663GAT_247_ngat), .B(G3768GAT_1363_ngat), .Y(G3836GAT_1398_gat) );
AND2XL U_g1368 (.A(G3764GAT_1364_ngat), .B(G3608GAT_1294_ngat), .Y(G3832GAT_1399_gat) );
AND2XL U_g1369 (.A(G615GAT_263_ngat), .B(G3764GAT_1364_ngat), .Y(G3831GAT_1400_gat) );
AND2XL U_g1370 (.A(G3760GAT_1365_ngat), .B(G3604GAT_1295_ngat), .Y(G3827GAT_1401_gat) );
AND2XL U_g1371 (.A(G567GAT_279_ngat), .B(G3760GAT_1365_ngat), .Y(G3826GAT_1402_gat) );
AND2XL U_g1372 (.A(G3894GAT_1367_ngat), .B(G3893GAT_1366_ngat), .Y(G3944GAT_1403_gat) );
AND2XL U_g1373 (.A(G3889GAT_1368_ngat), .B(G3818GAT_1345_ngat), .Y(G3942GAT_1404_gat) );
AND2XL U_g1374 (.A(G3815GAT_1346_ngat), .B(G3889GAT_1368_ngat), .Y(G3943GAT_1405_gat) );
AND2XL U_g1375 (.A(G3883GAT_1370_ngat), .B(G3886GAT_1369_ngat), .Y(G3938GAT_1406_gat) );
AND2XL U_g1376 (.A(G3882GAT_1380_ngat), .B(G3881GAT_1371_ngat), .Y(G3935GAT_1407_gat) );
AND2XL U_g1377 (.A(G3877GAT_1382_ngat), .B(G3693GAT_1299_ngat), .Y(G3932GAT_1408_gat) );
AND2XL U_g1378 (.A(G3877GAT_1382_ngat), .B(G3806GAT_1348_ngat), .Y(G3930GAT_1409_gat) );
AND2XL U_g1379 (.A(G3873GAT_1374_ngat), .B(G3872GAT_1373_ngat), .Y(G3923GAT_1410_gat) );
AND2XL U_g1380 (.A(G3868GAT_1375_ngat), .B(G3797GAT_1352_ngat), .Y(G3921GAT_1411_gat) );
AND2XL U_g1381 (.A(G3794GAT_1353_ngat), .B(G3868GAT_1375_ngat), .Y(G3922GAT_1412_gat) );
AND2XL U_g1382 (.A(G3862GAT_1386_ngat), .B(G3865GAT_1376_ngat), .Y(G3917GAT_1413_gat) );
AND2XL U_g1383 (.A(G3861GAT_1388_ngat), .B(G3860GAT_1377_ngat), .Y(G3914GAT_1414_gat) );
AND2XL U_g1384 (.A(G3856GAT_1390_ngat), .B(G3855GAT_1378_ngat), .Y(G3911GAT_1415_gat) );
AND2XL U_g1385 (.A(G3851GAT_1392_ngat), .B(G3850GAT_1379_ngat), .Y(G3908GAT_1416_gat) );
AND2XL U_g1386 (.A(G3846GAT_1394_ngat), .B(G3845GAT_1381_ngat), .Y(G3905GAT_1417_gat) );
AND2XL U_g1387 (.A(G1098GAT_102_ngat), .B(G3877GAT_1382_ngat), .Y(G3931GAT_1418_gat) );
AND2XL U_g1388 (.A(G3841GAT_1396_ngat), .B(G3840GAT_1383_ngat), .Y(G3902GAT_1419_gat) );
AND2XL U_g1389 (.A(G1050GAT_118_ngat), .B(G3874GAT_1372_ngat), .Y(G3926GAT_1420_gat) );
AND2XL U_g1390 (.A(G3836GAT_1398_ngat), .B(G3835GAT_1384_ngat), .Y(G3899GAT_1421_gat) );
AND2XL U_g1391 (.A(G3831GAT_1400_ngat), .B(G3830GAT_1385_ngat), .Y(G3896GAT_1422_gat) );
AND2XL U_g1392 (.A(G3826GAT_1402_ngat), .B(G3825GAT_1387_ngat), .Y(G3895GAT_1423_gat) );
AND2XL U_g1393 (.A(G3943GAT_1405_ngat), .B(G3942GAT_1404_ngat), .Y(G3998GAT_1424_gat) );
AND2XL U_g1394 (.A(G3938GAT_1406_ngat), .B(G3886GAT_1369_ngat), .Y(G3996GAT_1425_gat) );
AND2XL U_g1395 (.A(G3883GAT_1370_ngat), .B(G3938GAT_1406_ngat), .Y(G3997GAT_1426_gat) );
AND2XL U_g1396 (.A(G3932GAT_1408_ngat), .B(G3935GAT_1407_ngat), .Y(G3992GAT_1427_gat) );
AND2XL U_g1397 (.A(G3931GAT_1418_ngat), .B(G3930GAT_1409_ngat), .Y(G3989GAT_1428_gat) );
AND2XL U_g1398 (.A(G3926GAT_1420_ngat), .B(G3742GAT_1328_ngat), .Y(G3986GAT_1429_gat) );
AND2XL U_g1399 (.A(G3926GAT_1420_ngat), .B(G3874GAT_1372_ngat), .Y(G3984GAT_1430_gat) );
AND2XL U_g1400 (.A(G3922GAT_1412_ngat), .B(G3921GAT_1411_ngat), .Y(G3977GAT_1431_gat) );
AND2XL U_g1401 (.A(G3917GAT_1413_ngat), .B(G3865GAT_1376_ngat), .Y(G3975GAT_1432_gat) );
AND2XL U_g1402 (.A(G1245GAT_53_ngat), .B(G3944GAT_1403_ngat), .Y(G4001GAT_1433_gat) );
AND2XL U_g1403 (.A(G1050GAT_118_ngat), .B(G3926GAT_1420_ngat), .Y(G3985GAT_1434_gat) );
AND2XL U_g1404 (.A(G1002GAT_134_ngat), .B(G3923GAT_1410_ngat), .Y(G3980GAT_1435_gat) );
AND2XL U_g1405 (.A(G3862GAT_1386_ngat), .B(G3917GAT_1413_ngat), .Y(G3976GAT_1436_gat) );
AND2XL U_g1406 (.A(G3857GAT_1389_ngat), .B(G3914GAT_1414_ngat), .Y(G3971GAT_1437_gat) );
AND2XL U_g1407 (.A(G3852GAT_1391_ngat), .B(G3911GAT_1415_ngat), .Y(G3967GAT_1438_gat) );
AND2XL U_g1408 (.A(G3847GAT_1393_ngat), .B(G3908GAT_1416_ngat), .Y(G3963GAT_1439_gat) );
AND2XL U_g1409 (.A(G3842GAT_1395_ngat), .B(G3905GAT_1417_ngat), .Y(G3959GAT_1440_gat) );
AND2XL U_g1410 (.A(G3837GAT_1397_ngat), .B(G3902GAT_1419_ngat), .Y(G3955GAT_1441_gat) );
AND2XL U_g1411 (.A(G3832GAT_1399_ngat), .B(G3899GAT_1421_ngat), .Y(G3951GAT_1442_gat) );
AND2XL U_g1412 (.A(G3827GAT_1401_ngat), .B(G3896GAT_1422_ngat), .Y(G3947GAT_1443_gat) );
AND2XL U_g1413 (.A(G4001GAT_1433_ngat), .B(G3821GAT_1344_ngat), .Y(G4049GAT_1444_gat) );
AND2XL U_g1414 (.A(G4001GAT_1433_ngat), .B(G3944GAT_1403_ngat), .Y(G4047GAT_1445_gat) );
AND2XL U_g1415 (.A(G3997GAT_1426_ngat), .B(G3996GAT_1425_ngat), .Y(G4040GAT_1446_gat) );
AND2XL U_g1416 (.A(G3992GAT_1427_ngat), .B(G3935GAT_1407_ngat), .Y(G4038GAT_1447_gat) );
AND2XL U_g1417 (.A(G3932GAT_1408_ngat), .B(G3992GAT_1427_ngat), .Y(G4039GAT_1448_gat) );
AND2XL U_g1418 (.A(G3986GAT_1429_ngat), .B(G3989GAT_1428_ngat), .Y(G4034GAT_1449_gat) );
AND2XL U_g1419 (.A(G3985GAT_1434_ngat), .B(G3984GAT_1430_ngat), .Y(G4031GAT_1450_gat) );
AND2XL U_g1420 (.A(G3980GAT_1435_ngat), .B(G3800GAT_1351_ngat), .Y(G4028GAT_1451_gat) );
AND2XL U_g1421 (.A(G3980GAT_1435_ngat), .B(G3923GAT_1410_ngat), .Y(G4026GAT_1452_gat) );
AND2XL U_g1422 (.A(G3976GAT_1436_ngat), .B(G3975GAT_1432_ngat), .Y(G4019GAT_1453_gat) );
AND2XL U_g1423 (.A(G3971GAT_1437_ngat), .B(G3914GAT_1414_ngat), .Y(G4017GAT_1454_gat) );
AND2XL U_g1424 (.A(G1245GAT_53_ngat), .B(G4001GAT_1433_ngat), .Y(G4048GAT_1455_gat) );
AND2XL U_g1425 (.A(G3967GAT_1438_ngat), .B(G3911GAT_1415_ngat), .Y(G4015GAT_1456_gat) );
AND2XL U_g1426 (.A(G1197GAT_69_ngat), .B(G3998GAT_1424_ngat), .Y(G4043GAT_1457_gat) );
AND2XL U_g1427 (.A(G3963GAT_1439_ngat), .B(G3908GAT_1416_ngat), .Y(G4013GAT_1458_gat) );
AND2XL U_g1428 (.A(G3959GAT_1440_ngat), .B(G3905GAT_1417_ngat), .Y(G4011GAT_1459_gat) );
AND2XL U_g1429 (.A(G3955GAT_1441_ngat), .B(G3902GAT_1419_ngat), .Y(G4009GAT_1460_gat) );
AND2XL U_g1430 (.A(G3951GAT_1442_ngat), .B(G3899GAT_1421_ngat), .Y(G4007GAT_1461_gat) );
AND2XL U_g1431 (.A(G1002GAT_134_ngat), .B(G3980GAT_1435_ngat), .Y(G4027GAT_1462_gat) );
AND2XL U_g1432 (.A(G3947GAT_1443_ngat), .B(G3896GAT_1422_ngat), .Y(G4005GAT_1463_gat) );
AND2XL U_g1433 (.A(G954GAT_150_ngat), .B(G3977GAT_1431_ngat), .Y(G4022GAT_1464_gat) );
AND2XL U_g1434 (.A(G3857GAT_1389_ngat), .B(G3971GAT_1437_ngat), .Y(G4018GAT_1465_gat) );
AND2XL U_g1435 (.A(G3852GAT_1391_ngat), .B(G3967GAT_1438_ngat), .Y(G4016GAT_1466_gat) );
AND2XL U_g1436 (.A(G3847GAT_1393_ngat), .B(G3963GAT_1439_ngat), .Y(G4014GAT_1467_gat) );
AND2XL U_g1437 (.A(G3842GAT_1395_ngat), .B(G3959GAT_1440_ngat), .Y(G4012GAT_1468_gat) );
AND2XL U_g1438 (.A(G3837GAT_1397_ngat), .B(G3955GAT_1441_ngat), .Y(G4010GAT_1469_gat) );
AND2XL U_g1439 (.A(G3832GAT_1399_ngat), .B(G3951GAT_1442_ngat), .Y(G4008GAT_1470_gat) );
AND2XL U_g1440 (.A(G3827GAT_1401_ngat), .B(G3947GAT_1443_ngat), .Y(G4006GAT_1471_gat) );
AND2XL U_g1441 (.A(G4049GAT_1444_ngat), .B(G1293GAT_37_ngat), .Y(G4106GAT_1472_gat) );
AND2XL U_g1442 (.A(G4048GAT_1455_ngat), .B(G4047GAT_1445_ngat), .Y(G4103GAT_1473_gat) );
AND2XL U_g1443 (.A(G4043GAT_1457_ngat), .B(G3889GAT_1368_ngat), .Y(G4100GAT_1474_gat) );
AND2XL U_g1444 (.A(G4043GAT_1457_ngat), .B(G3998GAT_1424_ngat), .Y(G4098GAT_1475_gat) );
AND2XL U_g1445 (.A(G4039GAT_1448_ngat), .B(G4038GAT_1447_ngat), .Y(G4091GAT_1476_gat) );
AND2XL U_g1446 (.A(G4034GAT_1449_ngat), .B(G3989GAT_1428_ngat), .Y(G4089GAT_1477_gat) );
AND2XL U_g1447 (.A(G3986GAT_1429_ngat), .B(G4034GAT_1449_ngat), .Y(G4090GAT_1478_gat) );
AND2XL U_g1448 (.A(G4028GAT_1451_ngat), .B(G4031GAT_1450_ngat), .Y(G4085GAT_1479_gat) );
AND2XL U_g1449 (.A(G4027GAT_1462_ngat), .B(G4026GAT_1452_ngat), .Y(G4082GAT_1480_gat) );
AND2XL U_g1450 (.A(G4022GAT_1464_ngat), .B(G3868GAT_1375_ngat), .Y(G4079GAT_1481_gat) );
AND2XL U_g1451 (.A(G4022GAT_1464_ngat), .B(G3977GAT_1431_ngat), .Y(G4077GAT_1482_gat) );
AND2XL U_g1452 (.A(G4018GAT_1465_ngat), .B(G4017GAT_1454_ngat), .Y(G4070GAT_1483_gat) );
AND2XL U_g1453 (.A(G4016GAT_1466_ngat), .B(G4015GAT_1456_ngat), .Y(G4067GAT_1484_gat) );
AND2XL U_g1454 (.A(G1197GAT_69_ngat), .B(G4043GAT_1457_ngat), .Y(G4099GAT_1485_gat) );
AND2XL U_g1455 (.A(G4014GAT_1467_ngat), .B(G4013GAT_1458_ngat), .Y(G4064GAT_1486_gat) );
AND2XL U_g1456 (.A(G1149GAT_85_ngat), .B(G4040GAT_1446_ngat), .Y(G4094GAT_1487_gat) );
AND2XL U_g1457 (.A(G4012GAT_1468_ngat), .B(G4011GAT_1459_ngat), .Y(G4061GAT_1488_gat) );
AND2XL U_g1458 (.A(G4010GAT_1469_ngat), .B(G4009GAT_1460_ngat), .Y(G4058GAT_1489_gat) );
AND2XL U_g1459 (.A(G4008GAT_1470_ngat), .B(G4007GAT_1461_ngat), .Y(G4055GAT_1490_gat) );
AND2XL U_g1460 (.A(G4006GAT_1471_ngat), .B(G4005GAT_1463_ngat), .Y(G4052GAT_1491_gat) );
AND2XL U_g1461 (.A(G954GAT_150_ngat), .B(G4022GAT_1464_ngat), .Y(G4078GAT_1492_gat) );
AND2XL U_g1462 (.A(G906GAT_166_ngat), .B(G4019GAT_1453_ngat), .Y(G4073GAT_1493_gat) );
AND2XL U_g1463 (.A(G4106GAT_1472_ngat), .B(G1293GAT_37_ngat), .Y(G4171GAT_1494_gat) );
AND2XL U_g1464 (.A(G4049GAT_1444_ngat), .B(G4106GAT_1472_ngat), .Y(G4172GAT_1495_gat) );
AND2XL U_g1465 (.A(G4100GAT_1474_ngat), .B(G4103GAT_1473_ngat), .Y(G4167GAT_1496_gat) );
AND2XL U_g1466 (.A(G4099GAT_1485_ngat), .B(G4098GAT_1475_ngat), .Y(G4164GAT_1497_gat) );
AND2XL U_g1467 (.A(G4094GAT_1487_ngat), .B(G3938GAT_1406_ngat), .Y(G4161GAT_1498_gat) );
AND2XL U_g1468 (.A(G4094GAT_1487_ngat), .B(G4040GAT_1446_ngat), .Y(G4159GAT_1499_gat) );
AND2XL U_g1469 (.A(G4090GAT_1478_ngat), .B(G4089GAT_1477_ngat), .Y(G4152GAT_1500_gat) );
AND2XL U_g1470 (.A(G4085GAT_1479_ngat), .B(G4031GAT_1450_ngat), .Y(G4150GAT_1501_gat) );
AND2XL U_g1471 (.A(G4028GAT_1451_ngat), .B(G4085GAT_1479_ngat), .Y(G4151GAT_1502_gat) );
AND2XL U_g1472 (.A(G4079GAT_1481_ngat), .B(G4082GAT_1480_ngat), .Y(G4146GAT_1503_gat) );
AND2XL U_g1473 (.A(G4078GAT_1492_ngat), .B(G4077GAT_1482_ngat), .Y(G4143GAT_1504_gat) );
AND2XL U_g1474 (.A(G4073GAT_1493_ngat), .B(G3917GAT_1413_ngat), .Y(G4140GAT_1505_gat) );
AND2XL U_g1475 (.A(G4073GAT_1493_ngat), .B(G4019GAT_1453_ngat), .Y(G4138GAT_1506_gat) );
AND2XL U_g1476 (.A(G1149GAT_85_ngat), .B(G4094GAT_1487_ngat), .Y(G4160GAT_1507_gat) );
AND2XL U_g1477 (.A(G1101GAT_101_ngat), .B(G4091GAT_1476_ngat), .Y(G4155GAT_1508_gat) );
AND2XL U_g1478 (.A(G906GAT_166_ngat), .B(G4073GAT_1493_ngat), .Y(G4139GAT_1509_gat) );
AND2XL U_g1479 (.A(G858GAT_182_ngat), .B(G4070GAT_1483_ngat), .Y(G4134GAT_1510_gat) );
AND2XL U_g1480 (.A(G810GAT_198_ngat), .B(G4067GAT_1484_ngat), .Y(G4130GAT_1511_gat) );
AND2XL U_g1481 (.A(G762GAT_214_ngat), .B(G4064GAT_1486_ngat), .Y(G4126GAT_1512_gat) );
AND2XL U_g1482 (.A(G714GAT_230_ngat), .B(G4061GAT_1488_ngat), .Y(G4122GAT_1513_gat) );
AND2XL U_g1483 (.A(G666GAT_246_ngat), .B(G4058GAT_1489_ngat), .Y(G4118GAT_1514_gat) );
AND2XL U_g1484 (.A(G618GAT_262_ngat), .B(G4055GAT_1490_ngat), .Y(G4114GAT_1515_gat) );
AND2XL U_g1485 (.A(G570GAT_278_ngat), .B(G4052GAT_1491_ngat), .Y(G4110GAT_1516_gat) );
AND2XL U_g1486 (.A(G4172GAT_1495_ngat), .B(G4171GAT_1494_ngat), .Y(G4238GAT_1517_gat) );
AND2XL U_g1487 (.A(G4167GAT_1496_ngat), .B(G4103GAT_1473_ngat), .Y(G4236GAT_1518_gat) );
AND2XL U_g1488 (.A(G4100GAT_1474_ngat), .B(G4167GAT_1496_ngat), .Y(G4237GAT_1519_gat) );
AND2XL U_g1489 (.A(G4161GAT_1498_ngat), .B(G4164GAT_1497_ngat), .Y(G4232GAT_1520_gat) );
AND2XL U_g1490 (.A(G4160GAT_1507_ngat), .B(G4159GAT_1499_ngat), .Y(G4229GAT_1521_gat) );
AND2XL U_g1491 (.A(G4155GAT_1508_ngat), .B(G3992GAT_1427_ngat), .Y(G4226GAT_1522_gat) );
AND2XL U_g1492 (.A(G4155GAT_1508_ngat), .B(G4091GAT_1476_ngat), .Y(G4224GAT_1523_gat) );
AND2XL U_g1493 (.A(G4151GAT_1502_ngat), .B(G4150GAT_1501_ngat), .Y(G4217GAT_1524_gat) );
AND2XL U_g1494 (.A(G4146GAT_1503_ngat), .B(G4082GAT_1480_ngat), .Y(G4215GAT_1525_gat) );
AND2XL U_g1495 (.A(G4079GAT_1481_ngat), .B(G4146GAT_1503_ngat), .Y(G4216GAT_1526_gat) );
AND2XL U_g1496 (.A(G4140GAT_1505_ngat), .B(G4143GAT_1504_ngat), .Y(G4211GAT_1527_gat) );
AND2XL U_g1497 (.A(G4139GAT_1509_ngat), .B(G4138GAT_1506_ngat), .Y(G4208GAT_1528_gat) );
AND2XL U_g1498 (.A(G4134GAT_1510_ngat), .B(G4070GAT_1483_ngat), .Y(G4203GAT_1529_gat) );
AND2XL U_g1499 (.A(G4130GAT_1511_ngat), .B(G4067GAT_1484_ngat), .Y(G4198GAT_1530_gat) );
AND2XL U_g1500 (.A(G4126GAT_1512_ngat), .B(G4064GAT_1486_ngat), .Y(G4193GAT_1531_gat) );
AND2XL U_g1501 (.A(G4122GAT_1513_ngat), .B(G4061GAT_1488_ngat), .Y(G4188GAT_1532_gat) );
AND2XL U_g1502 (.A(G1101GAT_101_ngat), .B(G4155GAT_1508_ngat), .Y(G4225GAT_1533_gat) );
AND2XL U_g1503 (.A(G4118GAT_1514_ngat), .B(G4058GAT_1489_ngat), .Y(G4183GAT_1534_gat) );
AND2XL U_g1504 (.A(G1053GAT_117_ngat), .B(G4152GAT_1500_ngat), .Y(G4220GAT_1535_gat) );
AND2XL U_g1505 (.A(G4114GAT_1515_ngat), .B(G4055GAT_1490_ngat), .Y(G4178GAT_1536_gat) );
AND2XL U_g1506 (.A(G4110GAT_1516_ngat), .B(G4052GAT_1491_ngat), .Y(G4173GAT_1537_gat) );
AND2XL U_g1507 (.A(G4134GAT_1510_ngat), .B(G3971GAT_1437_ngat), .Y(G4205GAT_1538_gat) );
AND2XL U_g1508 (.A(G858GAT_182_ngat), .B(G4134GAT_1510_ngat), .Y(G4204GAT_1539_gat) );
AND2XL U_g1509 (.A(G4130GAT_1511_ngat), .B(G3967GAT_1438_ngat), .Y(G4200GAT_1540_gat) );
AND2XL U_g1510 (.A(G810GAT_198_ngat), .B(G4130GAT_1511_ngat), .Y(G4199GAT_1541_gat) );
AND2XL U_g1511 (.A(G4126GAT_1512_ngat), .B(G3963GAT_1439_ngat), .Y(G4195GAT_1542_gat) );
AND2XL U_g1512 (.A(G762GAT_214_ngat), .B(G4126GAT_1512_ngat), .Y(G4194GAT_1543_gat) );
AND2XL U_g1513 (.A(G4122GAT_1513_ngat), .B(G3959GAT_1440_ngat), .Y(G4190GAT_1544_gat) );
AND2XL U_g1514 (.A(G714GAT_230_ngat), .B(G4122GAT_1513_ngat), .Y(G4189GAT_1545_gat) );
AND2XL U_g1515 (.A(G4118GAT_1514_ngat), .B(G3955GAT_1441_ngat), .Y(G4185GAT_1546_gat) );
AND2XL U_g1516 (.A(G666GAT_246_ngat), .B(G4118GAT_1514_ngat), .Y(G4184GAT_1547_gat) );
AND2XL U_g1517 (.A(G4114GAT_1515_ngat), .B(G3951GAT_1442_ngat), .Y(G4180GAT_1548_gat) );
AND2XL U_g1518 (.A(G618GAT_262_ngat), .B(G4114GAT_1515_ngat), .Y(G4179GAT_1549_gat) );
AND2XL U_g1519 (.A(G4110GAT_1516_ngat), .B(G3947GAT_1443_ngat), .Y(G4175GAT_1550_gat) );
AND2XL U_g1520 (.A(G570GAT_278_ngat), .B(G4110GAT_1516_ngat), .Y(G4174GAT_1551_gat) );
AND2XL U_g1521 (.A(G4237GAT_1519_ngat), .B(G4236GAT_1518_ngat), .Y(G4287GAT_1552_gat) );
AND2XL U_g1522 (.A(G4232GAT_1520_ngat), .B(G4164GAT_1497_ngat), .Y(G4285GAT_1553_gat) );
AND2XL U_g1523 (.A(G4161GAT_1498_ngat), .B(G4232GAT_1520_ngat), .Y(G4286GAT_1554_gat) );
AND2XL U_g1524 (.A(G4226GAT_1522_ngat), .B(G4229GAT_1521_ngat), .Y(G4281GAT_1555_gat) );
AND2XL U_g1525 (.A(G4225GAT_1533_ngat), .B(G4224GAT_1523_ngat), .Y(G4278GAT_1556_gat) );
AND2XL U_g1526 (.A(G4220GAT_1535_ngat), .B(G4034GAT_1449_ngat), .Y(G4275GAT_1557_gat) );
AND2XL U_g1527 (.A(G4220GAT_1535_ngat), .B(G4152GAT_1500_ngat), .Y(G4273GAT_1558_gat) );
AND2XL U_g1528 (.A(G4216GAT_1526_ngat), .B(G4215GAT_1525_ngat), .Y(G4266GAT_1559_gat) );
AND2XL U_g1529 (.A(G4211GAT_1527_ngat), .B(G4143GAT_1504_ngat), .Y(G4264GAT_1560_gat) );
AND2XL U_g1530 (.A(G4140GAT_1505_ngat), .B(G4211GAT_1527_ngat), .Y(G4265GAT_1561_gat) );
AND2XL U_g1531 (.A(G4205GAT_1538_ngat), .B(G4208GAT_1528_ngat), .Y(G4260GAT_1562_gat) );
AND2XL U_g1532 (.A(G4204GAT_1539_ngat), .B(G4203GAT_1529_ngat), .Y(G4257GAT_1563_gat) );
AND2XL U_g1533 (.A(G1248GAT_52_ngat), .B(G4238GAT_1517_ngat), .Y(G4290GAT_1564_gat) );
AND2XL U_g1534 (.A(G4199GAT_1541_ngat), .B(G4198GAT_1530_ngat), .Y(G4254GAT_1565_gat) );
AND2XL U_g1535 (.A(G4194GAT_1543_ngat), .B(G4193GAT_1531_ngat), .Y(G4251GAT_1566_gat) );
AND2XL U_g1536 (.A(G4189GAT_1545_ngat), .B(G4188GAT_1532_ngat), .Y(G4248GAT_1567_gat) );
AND2XL U_g1537 (.A(G4184GAT_1547_ngat), .B(G4183GAT_1534_ngat), .Y(G4245GAT_1568_gat) );
AND2XL U_g1538 (.A(G1053GAT_117_ngat), .B(G4220GAT_1535_ngat), .Y(G4274GAT_1569_gat) );
AND2XL U_g1539 (.A(G4179GAT_1549_ngat), .B(G4178GAT_1536_ngat), .Y(G4242GAT_1570_gat) );
AND2XL U_g1540 (.A(G1005GAT_133_ngat), .B(G4217GAT_1524_ngat), .Y(G4269GAT_1571_gat) );
AND2XL U_g1541 (.A(G4174GAT_1551_ngat), .B(G4173GAT_1537_ngat), .Y(G4241GAT_1572_gat) );
AND2XL U_g1542 (.A(G4290GAT_1564_ngat), .B(G4106GAT_1472_ngat), .Y(G4350GAT_1573_gat) );
AND2XL U_g1543 (.A(G4290GAT_1564_ngat), .B(G4238GAT_1517_ngat), .Y(G4348GAT_1574_gat) );
AND2XL U_g1544 (.A(G4286GAT_1554_ngat), .B(G4285GAT_1553_ngat), .Y(G4341GAT_1575_gat) );
AND2XL U_g1545 (.A(G4281GAT_1555_ngat), .B(G4229GAT_1521_ngat), .Y(G4339GAT_1576_gat) );
AND2XL U_g1546 (.A(G4226GAT_1522_ngat), .B(G4281GAT_1555_ngat), .Y(G4340GAT_1577_gat) );
AND2XL U_g1547 (.A(G4275GAT_1557_ngat), .B(G4278GAT_1556_ngat), .Y(G4335GAT_1578_gat) );
AND2XL U_g1548 (.A(G4274GAT_1569_ngat), .B(G4273GAT_1558_ngat), .Y(G4332GAT_1579_gat) );
AND2XL U_g1549 (.A(G4269GAT_1571_ngat), .B(G4085GAT_1479_ngat), .Y(G4329GAT_1580_gat) );
AND2XL U_g1550 (.A(G4269GAT_1571_ngat), .B(G4217GAT_1524_ngat), .Y(G4327GAT_1581_gat) );
AND2XL U_g1551 (.A(G4265GAT_1561_ngat), .B(G4264GAT_1560_ngat), .Y(G4320GAT_1582_gat) );
AND2XL U_g1552 (.A(G4260GAT_1562_ngat), .B(G4208GAT_1528_ngat), .Y(G4318GAT_1583_gat) );
AND2XL U_g1553 (.A(G1248GAT_52_ngat), .B(G4290GAT_1564_ngat), .Y(G4349GAT_1584_gat) );
AND2XL U_g1554 (.A(G1200GAT_68_ngat), .B(G4287GAT_1552_ngat), .Y(G4344GAT_1585_gat) );
AND2XL U_g1555 (.A(G1005GAT_133_ngat), .B(G4269GAT_1571_ngat), .Y(G4328GAT_1586_gat) );
AND2XL U_g1556 (.A(G957GAT_149_ngat), .B(G4266GAT_1559_ngat), .Y(G4323GAT_1587_gat) );
AND2XL U_g1557 (.A(G4205GAT_1538_ngat), .B(G4260GAT_1562_ngat), .Y(G4319GAT_1588_gat) );
AND2XL U_g1558 (.A(G4200GAT_1540_ngat), .B(G4257GAT_1563_ngat), .Y(G4314GAT_1589_gat) );
AND2XL U_g1559 (.A(G4195GAT_1542_ngat), .B(G4254GAT_1565_ngat), .Y(G4310GAT_1590_gat) );
AND2XL U_g1560 (.A(G4190GAT_1544_ngat), .B(G4251GAT_1566_ngat), .Y(G4306GAT_1591_gat) );
AND2XL U_g1561 (.A(G4185GAT_1546_ngat), .B(G4248GAT_1567_ngat), .Y(G4302GAT_1592_gat) );
AND2XL U_g1562 (.A(G4180GAT_1548_ngat), .B(G4245GAT_1568_ngat), .Y(G4298GAT_1593_gat) );
AND2XL U_g1563 (.A(G4175GAT_1550_ngat), .B(G4242GAT_1570_ngat), .Y(G4294GAT_1594_gat) );
AND2XL U_g1564 (.A(G4350GAT_1573_ngat), .B(G1296GAT_36_ngat), .Y(G4401GAT_1595_gat) );
AND2XL U_g1565 (.A(G4349GAT_1584_ngat), .B(G4348GAT_1574_ngat), .Y(G4398GAT_1596_gat) );
AND2XL U_g1566 (.A(G4344GAT_1585_ngat), .B(G4167GAT_1496_ngat), .Y(G4395GAT_1597_gat) );
AND2XL U_g1567 (.A(G4344GAT_1585_ngat), .B(G4287GAT_1552_ngat), .Y(G4393GAT_1598_gat) );
AND2XL U_g1568 (.A(G4340GAT_1577_ngat), .B(G4339GAT_1576_ngat), .Y(G4386GAT_1599_gat) );
AND2XL U_g1569 (.A(G4335GAT_1578_ngat), .B(G4278GAT_1556_ngat), .Y(G4384GAT_1600_gat) );
AND2XL U_g1570 (.A(G4275GAT_1557_ngat), .B(G4335GAT_1578_ngat), .Y(G4385GAT_1601_gat) );
AND2XL U_g1571 (.A(G4329GAT_1580_ngat), .B(G4332GAT_1579_ngat), .Y(G4380GAT_1602_gat) );
AND2XL U_g1572 (.A(G4328GAT_1586_ngat), .B(G4327GAT_1581_ngat), .Y(G4377GAT_1603_gat) );
AND2XL U_g1573 (.A(G4323GAT_1587_ngat), .B(G4146GAT_1503_ngat), .Y(G4374GAT_1604_gat) );
AND2XL U_g1574 (.A(G4323GAT_1587_ngat), .B(G4266GAT_1559_ngat), .Y(G4372GAT_1605_gat) );
AND2XL U_g1575 (.A(G4319GAT_1588_ngat), .B(G4318GAT_1583_ngat), .Y(G4365GAT_1606_gat) );
AND2XL U_g1576 (.A(G4314GAT_1589_ngat), .B(G4257GAT_1563_ngat), .Y(G4363GAT_1607_gat) );
AND2XL U_g1577 (.A(G4310GAT_1590_ngat), .B(G4254GAT_1565_ngat), .Y(G4361GAT_1608_gat) );
AND2XL U_g1578 (.A(G1200GAT_68_ngat), .B(G4344GAT_1585_ngat), .Y(G4394GAT_1609_gat) );
AND2XL U_g1579 (.A(G4306GAT_1591_ngat), .B(G4251GAT_1566_ngat), .Y(G4359GAT_1610_gat) );
AND2XL U_g1580 (.A(G1152GAT_84_ngat), .B(G4341GAT_1575_ngat), .Y(G4389GAT_1611_gat) );
AND2XL U_g1581 (.A(G4302GAT_1592_ngat), .B(G4248GAT_1567_ngat), .Y(G4357GAT_1612_gat) );
AND2XL U_g1582 (.A(G4298GAT_1593_ngat), .B(G4245GAT_1568_ngat), .Y(G4355GAT_1613_gat) );
AND2XL U_g1583 (.A(G4294GAT_1594_ngat), .B(G4242GAT_1570_ngat), .Y(G4353GAT_1614_gat) );
AND2XL U_g1584 (.A(G957GAT_149_ngat), .B(G4323GAT_1587_ngat), .Y(G4373GAT_1615_gat) );
AND2XL U_g1585 (.A(G909GAT_165_ngat), .B(G4320GAT_1582_ngat), .Y(G4368GAT_1616_gat) );
AND2XL U_g1586 (.A(G4200GAT_1540_ngat), .B(G4314GAT_1589_ngat), .Y(G4364GAT_1617_gat) );
AND2XL U_g1587 (.A(G4195GAT_1542_ngat), .B(G4310GAT_1590_ngat), .Y(G4362GAT_1618_gat) );
AND2XL U_g1588 (.A(G4190GAT_1544_ngat), .B(G4306GAT_1591_ngat), .Y(G4360GAT_1619_gat) );
AND2XL U_g1589 (.A(G4185GAT_1546_ngat), .B(G4302GAT_1592_ngat), .Y(G4358GAT_1620_gat) );
AND2XL U_g1590 (.A(G4180GAT_1548_ngat), .B(G4298GAT_1593_ngat), .Y(G4356GAT_1621_gat) );
AND2XL U_g1591 (.A(G4175GAT_1550_ngat), .B(G4294GAT_1594_ngat), .Y(G4354GAT_1622_gat) );
AND2XL U_g1592 (.A(G4401GAT_1595_ngat), .B(G1296GAT_36_ngat), .Y(G4460GAT_1623_gat) );
AND2XL U_g1593 (.A(G4350GAT_1573_ngat), .B(G4401GAT_1595_ngat), .Y(G4461GAT_1624_gat) );
AND2XL U_g1594 (.A(G4395GAT_1597_ngat), .B(G4398GAT_1596_ngat), .Y(G4456GAT_1625_gat) );
AND2XL U_g1595 (.A(G4394GAT_1609_ngat), .B(G4393GAT_1598_ngat), .Y(G4453GAT_1626_gat) );
AND2XL U_g1596 (.A(G4389GAT_1611_ngat), .B(G4232GAT_1520_ngat), .Y(G4450GAT_1627_gat) );
AND2XL U_g1597 (.A(G4389GAT_1611_ngat), .B(G4341GAT_1575_ngat), .Y(G4448GAT_1628_gat) );
AND2XL U_g1598 (.A(G4385GAT_1601_ngat), .B(G4384GAT_1600_ngat), .Y(G4441GAT_1629_gat) );
AND2XL U_g1599 (.A(G4380GAT_1602_ngat), .B(G4332GAT_1579_ngat), .Y(G4439GAT_1630_gat) );
AND2XL U_g1600 (.A(G4329GAT_1580_ngat), .B(G4380GAT_1602_ngat), .Y(G4440GAT_1631_gat) );
AND2XL U_g1601 (.A(G4374GAT_1604_ngat), .B(G4377GAT_1603_ngat), .Y(G4435GAT_1632_gat) );
AND2XL U_g1602 (.A(G4373GAT_1615_ngat), .B(G4372GAT_1605_ngat), .Y(G4432GAT_1633_gat) );
AND2XL U_g1603 (.A(G4368GAT_1616_ngat), .B(G4211GAT_1527_ngat), .Y(G4429GAT_1634_gat) );
AND2XL U_g1604 (.A(G4368GAT_1616_ngat), .B(G4320GAT_1582_ngat), .Y(G4427GAT_1635_gat) );
AND2XL U_g1605 (.A(G4364GAT_1617_ngat), .B(G4363GAT_1607_ngat), .Y(G4420GAT_1636_gat) );
AND2XL U_g1606 (.A(G4362GAT_1618_ngat), .B(G4361GAT_1608_ngat), .Y(G4417GAT_1637_gat) );
AND2XL U_g1607 (.A(G4360GAT_1619_ngat), .B(G4359GAT_1610_ngat), .Y(G4414GAT_1638_gat) );
AND2XL U_g1608 (.A(G1152GAT_84_ngat), .B(G4389GAT_1611_ngat), .Y(G4449GAT_1639_gat) );
AND2XL U_g1609 (.A(G4358GAT_1620_ngat), .B(G4357GAT_1612_ngat), .Y(G4411GAT_1640_gat) );
AND2XL U_g1610 (.A(G1104GAT_100_ngat), .B(G4386GAT_1599_ngat), .Y(G4444GAT_1641_gat) );
AND2XL U_g1611 (.A(G4356GAT_1621_ngat), .B(G4355GAT_1613_ngat), .Y(G4408GAT_1642_gat) );
AND2XL U_g1612 (.A(G4354GAT_1622_ngat), .B(G4353GAT_1614_ngat), .Y(G4405GAT_1643_gat) );
AND2XL U_g1613 (.A(G909GAT_165_ngat), .B(G4368GAT_1616_ngat), .Y(G4428GAT_1644_gat) );
AND2XL U_g1614 (.A(G861GAT_181_ngat), .B(G4365GAT_1606_ngat), .Y(G4423GAT_1645_gat) );
AND2XL U_g1615 (.A(G4461GAT_1624_ngat), .B(G4460GAT_1623_ngat), .Y(G4521GAT_1646_gat) );
AND2XL U_g1616 (.A(G4456GAT_1625_ngat), .B(G4398GAT_1596_ngat), .Y(G4519GAT_1647_gat) );
AND2XL U_g1617 (.A(G4395GAT_1597_ngat), .B(G4456GAT_1625_ngat), .Y(G4520GAT_1648_gat) );
AND2XL U_g1618 (.A(G4450GAT_1627_ngat), .B(G4453GAT_1626_ngat), .Y(G4515GAT_1649_gat) );
AND2XL U_g1619 (.A(G4449GAT_1639_ngat), .B(G4448GAT_1628_ngat), .Y(G4512GAT_1650_gat) );
AND2XL U_g1620 (.A(G4444GAT_1641_ngat), .B(G4281GAT_1555_ngat), .Y(G4509GAT_1651_gat) );
AND2XL U_g1621 (.A(G4444GAT_1641_ngat), .B(G4386GAT_1599_ngat), .Y(G4507GAT_1652_gat) );
AND2XL U_g1622 (.A(G4440GAT_1631_ngat), .B(G4439GAT_1630_ngat), .Y(G4500GAT_1653_gat) );
AND2XL U_g1623 (.A(G4435GAT_1632_ngat), .B(G4377GAT_1603_ngat), .Y(G4498GAT_1654_gat) );
AND2XL U_g1624 (.A(G4374GAT_1604_ngat), .B(G4435GAT_1632_ngat), .Y(G4499GAT_1655_gat) );
AND2XL U_g1625 (.A(G4429GAT_1634_ngat), .B(G4432GAT_1633_ngat), .Y(G4494GAT_1656_gat) );
AND2XL U_g1626 (.A(G4428GAT_1644_ngat), .B(G4427GAT_1635_ngat), .Y(G4491GAT_1657_gat) );
AND2XL U_g1627 (.A(G4423GAT_1645_ngat), .B(G4260GAT_1562_ngat), .Y(G4488GAT_1658_gat) );
AND2XL U_g1628 (.A(G4423GAT_1645_ngat), .B(G4365GAT_1606_ngat), .Y(G4486GAT_1659_gat) );
AND2XL U_g1629 (.A(G1104GAT_100_ngat), .B(G4444GAT_1641_ngat), .Y(G4508GAT_1660_gat) );
AND2XL U_g1630 (.A(G1056GAT_116_ngat), .B(G4441GAT_1629_ngat), .Y(G4503GAT_1661_gat) );
AND2XL U_g1631 (.A(G861GAT_181_ngat), .B(G4423GAT_1645_ngat), .Y(G4487GAT_1662_gat) );
AND2XL U_g1632 (.A(G813GAT_197_ngat), .B(G4420GAT_1636_ngat), .Y(G4482GAT_1663_gat) );
AND2XL U_g1633 (.A(G765GAT_213_ngat), .B(G4417GAT_1637_ngat), .Y(G4478GAT_1664_gat) );
AND2XL U_g1634 (.A(G717GAT_229_ngat), .B(G4414GAT_1638_ngat), .Y(G4474GAT_1665_gat) );
AND2XL U_g1635 (.A(G669GAT_245_ngat), .B(G4411GAT_1640_ngat), .Y(G4470GAT_1666_gat) );
AND2XL U_g1636 (.A(G621GAT_261_ngat), .B(G4408GAT_1642_ngat), .Y(G4466GAT_1667_gat) );
AND2XL U_g1637 (.A(G573GAT_277_ngat), .B(G4405GAT_1643_ngat), .Y(G4462GAT_1668_gat) );
AND2XL U_g1638 (.A(G4520GAT_1648_ngat), .B(G4519GAT_1647_ngat), .Y(G4584GAT_1669_gat) );
AND2XL U_g1639 (.A(G4515GAT_1649_ngat), .B(G4453GAT_1626_ngat), .Y(G4582GAT_1670_gat) );
AND2XL U_g1640 (.A(G4450GAT_1627_ngat), .B(G4515GAT_1649_ngat), .Y(G4583GAT_1671_gat) );
AND2XL U_g1641 (.A(G4509GAT_1651_ngat), .B(G4512GAT_1650_ngat), .Y(G4578GAT_1672_gat) );
AND2XL U_g1642 (.A(G4508GAT_1660_ngat), .B(G4507GAT_1652_ngat), .Y(G4575GAT_1673_gat) );
AND2XL U_g1643 (.A(G4503GAT_1661_ngat), .B(G4335GAT_1578_ngat), .Y(G4572GAT_1674_gat) );
AND2XL U_g1644 (.A(G4503GAT_1661_ngat), .B(G4441GAT_1629_ngat), .Y(G4570GAT_1675_gat) );
AND2XL U_g1645 (.A(G4499GAT_1655_ngat), .B(G4498GAT_1654_ngat), .Y(G4563GAT_1676_gat) );
AND2XL U_g1646 (.A(G4494GAT_1656_ngat), .B(G4432GAT_1633_ngat), .Y(G4561GAT_1677_gat) );
AND2XL U_g1647 (.A(G4429GAT_1634_ngat), .B(G4494GAT_1656_ngat), .Y(G4562GAT_1678_gat) );
AND2XL U_g1648 (.A(G4488GAT_1658_ngat), .B(G4491GAT_1657_ngat), .Y(G4557GAT_1679_gat) );
AND2XL U_g1649 (.A(G4487GAT_1662_ngat), .B(G4486GAT_1659_ngat), .Y(G4554GAT_1680_gat) );
AND2XL U_g1650 (.A(G4482GAT_1663_ngat), .B(G4420GAT_1636_ngat), .Y(G4549GAT_1681_gat) );
AND2XL U_g1651 (.A(G1251GAT_51_ngat), .B(G4521GAT_1646_ngat), .Y(G4587GAT_1682_gat) );
AND2XL U_g1652 (.A(G4478GAT_1664_ngat), .B(G4417GAT_1637_ngat), .Y(G4544GAT_1683_gat) );
AND2XL U_g1653 (.A(G4474GAT_1665_ngat), .B(G4414GAT_1638_ngat), .Y(G4539GAT_1684_gat) );
AND2XL U_g1654 (.A(G4470GAT_1666_ngat), .B(G4411GAT_1640_ngat), .Y(G4534GAT_1685_gat) );
AND2XL U_g1655 (.A(G4466GAT_1667_ngat), .B(G4408GAT_1642_ngat), .Y(G4529GAT_1686_gat) );
AND2XL U_g1656 (.A(G1056GAT_116_ngat), .B(G4503GAT_1661_ngat), .Y(G4571GAT_1687_gat) );
AND2XL U_g1657 (.A(G4462GAT_1668_ngat), .B(G4405GAT_1643_ngat), .Y(G4524GAT_1688_gat) );
AND2XL U_g1658 (.A(G1008GAT_132_ngat), .B(G4500GAT_1653_ngat), .Y(G4566GAT_1689_gat) );
AND2XL U_g1659 (.A(G4482GAT_1663_ngat), .B(G4314GAT_1589_ngat), .Y(G4551GAT_1690_gat) );
AND2XL U_g1660 (.A(G813GAT_197_ngat), .B(G4482GAT_1663_ngat), .Y(G4550GAT_1691_gat) );
AND2XL U_g1661 (.A(G4478GAT_1664_ngat), .B(G4310GAT_1590_ngat), .Y(G4546GAT_1692_gat) );
AND2XL U_g1662 (.A(G765GAT_213_ngat), .B(G4478GAT_1664_ngat), .Y(G4545GAT_1693_gat) );
AND2XL U_g1663 (.A(G4474GAT_1665_ngat), .B(G4306GAT_1591_ngat), .Y(G4541GAT_1694_gat) );
AND2XL U_g1664 (.A(G717GAT_229_ngat), .B(G4474GAT_1665_ngat), .Y(G4540GAT_1695_gat) );
AND2XL U_g1665 (.A(G4470GAT_1666_ngat), .B(G4302GAT_1592_ngat), .Y(G4536GAT_1696_gat) );
AND2XL U_g1666 (.A(G669GAT_245_ngat), .B(G4470GAT_1666_ngat), .Y(G4535GAT_1697_gat) );
AND2XL U_g1667 (.A(G4466GAT_1667_ngat), .B(G4298GAT_1593_ngat), .Y(G4531GAT_1698_gat) );
AND2XL U_g1668 (.A(G621GAT_261_ngat), .B(G4466GAT_1667_ngat), .Y(G4530GAT_1699_gat) );
AND2XL U_g1669 (.A(G4462GAT_1668_ngat), .B(G4294GAT_1594_ngat), .Y(G4526GAT_1700_gat) );
AND2XL U_g1670 (.A(G573GAT_277_ngat), .B(G4462GAT_1668_ngat), .Y(G4525GAT_1701_gat) );
AND2XL U_g1671 (.A(G4587GAT_1682_ngat), .B(G4401GAT_1595_ngat), .Y(G4643GAT_1702_gat) );
AND2XL U_g1672 (.A(G4587GAT_1682_ngat), .B(G4521GAT_1646_ngat), .Y(G4641GAT_1703_gat) );
AND2XL U_g1673 (.A(G4583GAT_1671_ngat), .B(G4582GAT_1670_ngat), .Y(G4634GAT_1704_gat) );
AND2XL U_g1674 (.A(G4578GAT_1672_ngat), .B(G4512GAT_1650_ngat), .Y(G4632GAT_1705_gat) );
AND2XL U_g1675 (.A(G4509GAT_1651_ngat), .B(G4578GAT_1672_ngat), .Y(G4633GAT_1706_gat) );
AND2XL U_g1676 (.A(G4572GAT_1674_ngat), .B(G4575GAT_1673_ngat), .Y(G4628GAT_1707_gat) );
AND2XL U_g1677 (.A(G4571GAT_1687_ngat), .B(G4570GAT_1675_ngat), .Y(G4625GAT_1708_gat) );
AND2XL U_g1678 (.A(G4566GAT_1689_ngat), .B(G4380GAT_1602_ngat), .Y(G4622GAT_1709_gat) );
AND2XL U_g1679 (.A(G4566GAT_1689_ngat), .B(G4500GAT_1653_ngat), .Y(G4620GAT_1710_gat) );
AND2XL U_g1680 (.A(G4562GAT_1678_ngat), .B(G4561GAT_1677_ngat), .Y(G4613GAT_1711_gat) );
AND2XL U_g1681 (.A(G4557GAT_1679_ngat), .B(G4491GAT_1657_ngat), .Y(G4611GAT_1712_gat) );
AND2XL U_g1682 (.A(G4488GAT_1658_ngat), .B(G4557GAT_1679_ngat), .Y(G4612GAT_1713_gat) );
AND2XL U_g1683 (.A(G4551GAT_1690_ngat), .B(G4554GAT_1680_ngat), .Y(G4607GAT_1714_gat) );
AND2XL U_g1684 (.A(G4550GAT_1691_ngat), .B(G4549GAT_1681_ngat), .Y(G4604GAT_1715_gat) );
AND2XL U_g1685 (.A(G1251GAT_51_ngat), .B(G4587GAT_1682_ngat), .Y(G4642GAT_1716_gat) );
AND2XL U_g1686 (.A(G4545GAT_1693_ngat), .B(G4544GAT_1683_ngat), .Y(G4601GAT_1717_gat) );
AND2XL U_g1687 (.A(G1203GAT_67_ngat), .B(G4584GAT_1669_ngat), .Y(G4637GAT_1718_gat) );
AND2XL U_g1688 (.A(G4540GAT_1695_ngat), .B(G4539GAT_1684_ngat), .Y(G4598GAT_1719_gat) );
AND2XL U_g1689 (.A(G4535GAT_1697_ngat), .B(G4534GAT_1685_ngat), .Y(G4595GAT_1720_gat) );
AND2XL U_g1690 (.A(G4530GAT_1699_ngat), .B(G4529GAT_1686_ngat), .Y(G4592GAT_1721_gat) );
AND2XL U_g1691 (.A(G4525GAT_1701_ngat), .B(G4524GAT_1688_ngat), .Y(G4591GAT_1722_gat) );
AND2XL U_g1692 (.A(G1008GAT_132_ngat), .B(G4566GAT_1689_ngat), .Y(G4621GAT_1723_gat) );
AND2XL U_g1693 (.A(G960GAT_148_ngat), .B(G4563GAT_1676_ngat), .Y(G4616GAT_1724_gat) );
AND2XL U_g1694 (.A(G4643GAT_1702_ngat), .B(G1299GAT_35_ngat), .Y(G4704GAT_1725_gat) );
AND2XL U_g1695 (.A(G4642GAT_1716_ngat), .B(G4641GAT_1703_ngat), .Y(G4701GAT_1726_gat) );
AND2XL U_g1696 (.A(G4637GAT_1718_ngat), .B(G4456GAT_1625_ngat), .Y(G4698GAT_1727_gat) );
AND2XL U_g1697 (.A(G4637GAT_1718_ngat), .B(G4584GAT_1669_ngat), .Y(G4696GAT_1728_gat) );
AND2XL U_g1698 (.A(G4633GAT_1706_ngat), .B(G4632GAT_1705_ngat), .Y(G4689GAT_1729_gat) );
AND2XL U_g1699 (.A(G4628GAT_1707_ngat), .B(G4575GAT_1673_ngat), .Y(G4687GAT_1730_gat) );
AND2XL U_g1700 (.A(G4572GAT_1674_ngat), .B(G4628GAT_1707_ngat), .Y(G4688GAT_1731_gat) );
AND2XL U_g1701 (.A(G4622GAT_1709_ngat), .B(G4625GAT_1708_ngat), .Y(G4683GAT_1732_gat) );
AND2XL U_g1702 (.A(G4621GAT_1723_ngat), .B(G4620GAT_1710_ngat), .Y(G4680GAT_1733_gat) );
AND2XL U_g1703 (.A(G4616GAT_1724_ngat), .B(G4435GAT_1632_ngat), .Y(G4677GAT_1734_gat) );
AND2XL U_g1704 (.A(G4616GAT_1724_ngat), .B(G4563GAT_1676_ngat), .Y(G4675GAT_1735_gat) );
AND2XL U_g1705 (.A(G4612GAT_1713_ngat), .B(G4611GAT_1712_ngat), .Y(G4668GAT_1736_gat) );
AND2XL U_g1706 (.A(G4607GAT_1714_ngat), .B(G4554GAT_1680_ngat), .Y(G4666GAT_1737_gat) );
AND2XL U_g1707 (.A(G1203GAT_67_ngat), .B(G4637GAT_1718_ngat), .Y(G4697GAT_1738_gat) );
AND2XL U_g1708 (.A(G1155GAT_83_ngat), .B(G4634GAT_1704_ngat), .Y(G4692GAT_1739_gat) );
AND2XL U_g1709 (.A(G960GAT_148_ngat), .B(G4616GAT_1724_ngat), .Y(G4676GAT_1740_gat) );
AND2XL U_g1710 (.A(G912GAT_164_ngat), .B(G4613GAT_1711_ngat), .Y(G4671GAT_1741_gat) );
AND2XL U_g1711 (.A(G4551GAT_1690_ngat), .B(G4607GAT_1714_ngat), .Y(G4667GAT_1742_gat) );
AND2XL U_g1712 (.A(G4546GAT_1692_ngat), .B(G4604GAT_1715_ngat), .Y(G4662GAT_1743_gat) );
AND2XL U_g1713 (.A(G4541GAT_1694_ngat), .B(G4601GAT_1717_ngat), .Y(G4658GAT_1744_gat) );
AND2XL U_g1714 (.A(G4536GAT_1696_ngat), .B(G4598GAT_1719_ngat), .Y(G4654GAT_1745_gat) );
AND2XL U_g1715 (.A(G4531GAT_1698_ngat), .B(G4595GAT_1720_ngat), .Y(G4650GAT_1746_gat) );
AND2XL U_g1716 (.A(G4526GAT_1700_ngat), .B(G4592GAT_1721_ngat), .Y(G4646GAT_1747_gat) );
AND2XL U_g1717 (.A(G4704GAT_1725_ngat), .B(G1299GAT_35_ngat), .Y(G4758GAT_1748_gat) );
AND2XL U_g1718 (.A(G4643GAT_1702_ngat), .B(G4704GAT_1725_ngat), .Y(G4759GAT_1749_gat) );
AND2XL U_g1719 (.A(G4698GAT_1727_ngat), .B(G4701GAT_1726_ngat), .Y(G4754GAT_1750_gat) );
AND2XL U_g1720 (.A(G4697GAT_1738_ngat), .B(G4696GAT_1728_ngat), .Y(G4751GAT_1751_gat) );
AND2XL U_g1721 (.A(G4692GAT_1739_ngat), .B(G4515GAT_1649_ngat), .Y(G4748GAT_1752_gat) );
AND2XL U_g1722 (.A(G4692GAT_1739_ngat), .B(G4634GAT_1704_ngat), .Y(G4746GAT_1753_gat) );
AND2XL U_g1723 (.A(G4688GAT_1731_ngat), .B(G4687GAT_1730_ngat), .Y(G4739GAT_1754_gat) );
AND2XL U_g1724 (.A(G4683GAT_1732_ngat), .B(G4625GAT_1708_ngat), .Y(G4737GAT_1755_gat) );
AND2XL U_g1725 (.A(G4622GAT_1709_ngat), .B(G4683GAT_1732_ngat), .Y(G4738GAT_1756_gat) );
AND2XL U_g1726 (.A(G4677GAT_1734_ngat), .B(G4680GAT_1733_ngat), .Y(G4733GAT_1757_gat) );
AND2XL U_g1727 (.A(G4676GAT_1740_ngat), .B(G4675GAT_1735_ngat), .Y(G4730GAT_1758_gat) );
AND2XL U_g1728 (.A(G4671GAT_1741_ngat), .B(G4494GAT_1656_ngat), .Y(G4727GAT_1759_gat) );
AND2XL U_g1729 (.A(G4671GAT_1741_ngat), .B(G4613GAT_1711_ngat), .Y(G4725GAT_1760_gat) );
AND2XL U_g1730 (.A(G4667GAT_1742_ngat), .B(G4666GAT_1737_ngat), .Y(G4718GAT_1761_gat) );
AND2XL U_g1731 (.A(G4662GAT_1743_ngat), .B(G4604GAT_1715_ngat), .Y(G4716GAT_1762_gat) );
AND2XL U_g1732 (.A(G4658GAT_1744_ngat), .B(G4601GAT_1717_ngat), .Y(G4714GAT_1763_gat) );
AND2XL U_g1733 (.A(G4654GAT_1745_ngat), .B(G4598GAT_1719_ngat), .Y(G4712GAT_1764_gat) );
AND2XL U_g1734 (.A(G1155GAT_83_ngat), .B(G4692GAT_1739_ngat), .Y(G4747GAT_1765_gat) );
AND2XL U_g1735 (.A(G4650GAT_1746_ngat), .B(G4595GAT_1720_ngat), .Y(G4710GAT_1766_gat) );
AND2XL U_g1736 (.A(G1107GAT_99_ngat), .B(G4689GAT_1729_ngat), .Y(G4742GAT_1767_gat) );
AND2XL U_g1737 (.A(G4646GAT_1747_ngat), .B(G4592GAT_1721_ngat), .Y(G4708GAT_1768_gat) );
AND2XL U_g1738 (.A(G912GAT_164_ngat), .B(G4671GAT_1741_ngat), .Y(G4726GAT_1769_gat) );
AND2XL U_g1739 (.A(G864GAT_180_ngat), .B(G4668GAT_1736_ngat), .Y(G4721GAT_1770_gat) );
AND2XL U_g1740 (.A(G4546GAT_1692_ngat), .B(G4662GAT_1743_ngat), .Y(G4717GAT_1771_gat) );
AND2XL U_g1741 (.A(G4541GAT_1694_ngat), .B(G4658GAT_1744_ngat), .Y(G4715GAT_1772_gat) );
AND2XL U_g1742 (.A(G4536GAT_1696_ngat), .B(G4654GAT_1745_ngat), .Y(G4713GAT_1773_gat) );
AND2XL U_g1743 (.A(G4531GAT_1698_ngat), .B(G4650GAT_1746_ngat), .Y(G4711GAT_1774_gat) );
AND2XL U_g1744 (.A(G4526GAT_1700_ngat), .B(G4646GAT_1747_ngat), .Y(G4709GAT_1775_gat) );
AND2XL U_g1745 (.A(G4759GAT_1749_ngat), .B(G4758GAT_1748_ngat), .Y(G4814GAT_1776_gat) );
AND2XL U_g1746 (.A(G4754GAT_1750_ngat), .B(G4701GAT_1726_ngat), .Y(G4812GAT_1777_gat) );
AND2XL U_g1747 (.A(G4698GAT_1727_ngat), .B(G4754GAT_1750_ngat), .Y(G4813GAT_1778_gat) );
AND2XL U_g1748 (.A(G4748GAT_1752_ngat), .B(G4751GAT_1751_ngat), .Y(G4808GAT_1779_gat) );
AND2XL U_g1749 (.A(G4747GAT_1765_ngat), .B(G4746GAT_1753_ngat), .Y(G4805GAT_1780_gat) );
AND2XL U_g1750 (.A(G4742GAT_1767_ngat), .B(G4578GAT_1672_ngat), .Y(G4802GAT_1781_gat) );
AND2XL U_g1751 (.A(G4742GAT_1767_ngat), .B(G4689GAT_1729_ngat), .Y(G4800GAT_1782_gat) );
AND2XL U_g1752 (.A(G4738GAT_1756_ngat), .B(G4737GAT_1755_ngat), .Y(G4793GAT_1783_gat) );
AND2XL U_g1753 (.A(G4733GAT_1757_ngat), .B(G4680GAT_1733_ngat), .Y(G4791GAT_1784_gat) );
AND2XL U_g1754 (.A(G4677GAT_1734_ngat), .B(G4733GAT_1757_ngat), .Y(G4792GAT_1785_gat) );
AND2XL U_g1755 (.A(G4727GAT_1759_ngat), .B(G4730GAT_1758_ngat), .Y(G4787GAT_1786_gat) );
AND2XL U_g1756 (.A(G4726GAT_1769_ngat), .B(G4725GAT_1760_ngat), .Y(G4784GAT_1787_gat) );
AND2XL U_g1757 (.A(G4721GAT_1770_ngat), .B(G4557GAT_1679_ngat), .Y(G4781GAT_1788_gat) );
AND2XL U_g1758 (.A(G4721GAT_1770_ngat), .B(G4668GAT_1736_ngat), .Y(G4779GAT_1789_gat) );
AND2XL U_g1759 (.A(G4717GAT_1771_ngat), .B(G4716GAT_1762_ngat), .Y(G4772GAT_1790_gat) );
AND2XL U_g1760 (.A(G4715GAT_1772_ngat), .B(G4714GAT_1763_ngat), .Y(G4769GAT_1791_gat) );
AND2XL U_g1761 (.A(G4713GAT_1773_ngat), .B(G4712GAT_1764_ngat), .Y(G4766GAT_1792_gat) );
AND2XL U_g1762 (.A(G4711GAT_1774_ngat), .B(G4710GAT_1766_ngat), .Y(G4763GAT_1793_gat) );
AND2XL U_g1763 (.A(G1107GAT_99_ngat), .B(G4742GAT_1767_ngat), .Y(G4801GAT_1794_gat) );
AND2XL U_g1764 (.A(G4709GAT_1775_ngat), .B(G4708GAT_1768_ngat), .Y(G4760GAT_1795_gat) );
AND2XL U_g1765 (.A(G1059GAT_115_ngat), .B(G4739GAT_1754_ngat), .Y(G4796GAT_1796_gat) );
AND2XL U_g1766 (.A(G864GAT_180_ngat), .B(G4721GAT_1770_ngat), .Y(G4780GAT_1797_gat) );
AND2XL U_g1767 (.A(G816GAT_196_ngat), .B(G4718GAT_1761_ngat), .Y(G4775GAT_1798_gat) );
AND2XL U_g1768 (.A(G4813GAT_1778_ngat), .B(G4812GAT_1777_ngat), .Y(G4872GAT_1799_gat) );
AND2XL U_g1769 (.A(G4808GAT_1779_ngat), .B(G4751GAT_1751_ngat), .Y(G4870GAT_1800_gat) );
AND2XL U_g1770 (.A(G4748GAT_1752_ngat), .B(G4808GAT_1779_ngat), .Y(G4871GAT_1801_gat) );
AND2XL U_g1771 (.A(G4802GAT_1781_ngat), .B(G4805GAT_1780_ngat), .Y(G4866GAT_1802_gat) );
AND2XL U_g1772 (.A(G4801GAT_1794_ngat), .B(G4800GAT_1782_ngat), .Y(G4863GAT_1803_gat) );
AND2XL U_g1773 (.A(G4796GAT_1796_ngat), .B(G4628GAT_1707_ngat), .Y(G4860GAT_1804_gat) );
AND2XL U_g1774 (.A(G4796GAT_1796_ngat), .B(G4739GAT_1754_ngat), .Y(G4858GAT_1805_gat) );
AND2XL U_g1775 (.A(G4792GAT_1785_ngat), .B(G4791GAT_1784_ngat), .Y(G4851GAT_1806_gat) );
AND2XL U_g1776 (.A(G4787GAT_1786_ngat), .B(G4730GAT_1758_ngat), .Y(G4849GAT_1807_gat) );
AND2XL U_g1777 (.A(G4727GAT_1759_ngat), .B(G4787GAT_1786_ngat), .Y(G4850GAT_1808_gat) );
AND2XL U_g1778 (.A(G4781GAT_1788_ngat), .B(G4784GAT_1787_ngat), .Y(G4845GAT_1809_gat) );
AND2XL U_g1779 (.A(G4780GAT_1797_ngat), .B(G4779GAT_1789_ngat), .Y(G4842GAT_1810_gat) );
AND2XL U_g1780 (.A(G4775GAT_1798_ngat), .B(G4607GAT_1714_ngat), .Y(G4839GAT_1811_gat) );
AND2XL U_g1781 (.A(G4775GAT_1798_ngat), .B(G4718GAT_1761_ngat), .Y(G4837GAT_1812_gat) );
AND2XL U_g1782 (.A(G1254GAT_50_ngat), .B(G4814GAT_1776_ngat), .Y(G4875GAT_1813_gat) );
AND2XL U_g1783 (.A(G1059GAT_115_ngat), .B(G4796GAT_1796_ngat), .Y(G4859GAT_1814_gat) );
AND2XL U_g1784 (.A(G1011GAT_131_ngat), .B(G4793GAT_1783_ngat), .Y(G4854GAT_1815_gat) );
AND2XL U_g1785 (.A(G816GAT_196_ngat), .B(G4775GAT_1798_ngat), .Y(G4838GAT_1816_gat) );
AND2XL U_g1786 (.A(G768GAT_212_ngat), .B(G4772GAT_1790_ngat), .Y(G4833GAT_1817_gat) );
AND2XL U_g1787 (.A(G720GAT_228_ngat), .B(G4769GAT_1791_ngat), .Y(G4829GAT_1818_gat) );
AND2XL U_g1788 (.A(G672GAT_244_ngat), .B(G4766GAT_1792_ngat), .Y(G4825GAT_1819_gat) );
AND2XL U_g1789 (.A(G624GAT_260_ngat), .B(G4763GAT_1793_ngat), .Y(G4821GAT_1820_gat) );
AND2XL U_g1790 (.A(G576GAT_276_ngat), .B(G4760GAT_1795_ngat), .Y(G4817GAT_1821_gat) );
AND2XL U_g1791 (.A(G4875GAT_1813_ngat), .B(G4704GAT_1725_ngat), .Y(G4943GAT_1822_gat) );
AND2XL U_g1792 (.A(G4875GAT_1813_ngat), .B(G4814GAT_1776_ngat), .Y(G4941GAT_1823_gat) );
AND2XL U_g1793 (.A(G4871GAT_1801_ngat), .B(G4870GAT_1800_ngat), .Y(G4934GAT_1824_gat) );
AND2XL U_g1794 (.A(G4866GAT_1802_ngat), .B(G4805GAT_1780_ngat), .Y(G4932GAT_1825_gat) );
AND2XL U_g1795 (.A(G4802GAT_1781_ngat), .B(G4866GAT_1802_ngat), .Y(G4933GAT_1826_gat) );
AND2XL U_g1796 (.A(G4860GAT_1804_ngat), .B(G4863GAT_1803_ngat), .Y(G4928GAT_1827_gat) );
AND2XL U_g1797 (.A(G4859GAT_1814_ngat), .B(G4858GAT_1805_ngat), .Y(G4925GAT_1828_gat) );
AND2XL U_g1798 (.A(G4854GAT_1815_ngat), .B(G4683GAT_1732_ngat), .Y(G4922GAT_1829_gat) );
AND2XL U_g1799 (.A(G4854GAT_1815_ngat), .B(G4793GAT_1783_ngat), .Y(G4920GAT_1830_gat) );
AND2XL U_g1800 (.A(G4850GAT_1808_ngat), .B(G4849GAT_1807_ngat), .Y(G4913GAT_1831_gat) );
AND2XL U_g1801 (.A(G4845GAT_1809_ngat), .B(G4784GAT_1787_ngat), .Y(G4911GAT_1832_gat) );
AND2XL U_g1802 (.A(G4781GAT_1788_ngat), .B(G4845GAT_1809_ngat), .Y(G4912GAT_1833_gat) );
AND2XL U_g1803 (.A(G4839GAT_1811_ngat), .B(G4842GAT_1810_ngat), .Y(G4907GAT_1834_gat) );
AND2XL U_g1804 (.A(G4838GAT_1816_ngat), .B(G4837GAT_1812_ngat), .Y(G4904GAT_1835_gat) );
AND2XL U_g1805 (.A(G4833GAT_1817_ngat), .B(G4772GAT_1790_ngat), .Y(G4899GAT_1836_gat) );
AND2XL U_g1806 (.A(G1254GAT_50_ngat), .B(G4875GAT_1813_ngat), .Y(G4942GAT_1837_gat) );
AND2XL U_g1807 (.A(G4829GAT_1818_ngat), .B(G4769GAT_1791_ngat), .Y(G4894GAT_1838_gat) );
AND2XL U_g1808 (.A(G1206GAT_66_ngat), .B(G4872GAT_1799_ngat), .Y(G4937GAT_1839_gat) );
AND2XL U_g1809 (.A(G4825GAT_1819_ngat), .B(G4766GAT_1792_ngat), .Y(G4889GAT_1840_gat) );
AND2XL U_g1810 (.A(G4821GAT_1820_ngat), .B(G4763GAT_1793_ngat), .Y(G4884GAT_1841_gat) );
AND2XL U_g1811 (.A(G4817GAT_1821_ngat), .B(G4760GAT_1795_ngat), .Y(G4879GAT_1842_gat) );
AND2XL U_g1812 (.A(G1011GAT_131_ngat), .B(G4854GAT_1815_ngat), .Y(G4921GAT_1843_gat) );
AND2XL U_g1813 (.A(G963GAT_147_ngat), .B(G4851GAT_1806_ngat), .Y(G4916GAT_1844_gat) );
AND2XL U_g1814 (.A(G4833GAT_1817_ngat), .B(G4662GAT_1743_ngat), .Y(G4901GAT_1845_gat) );
AND2XL U_g1815 (.A(G768GAT_212_ngat), .B(G4833GAT_1817_ngat), .Y(G4900GAT_1846_gat) );
AND2XL U_g1816 (.A(G4829GAT_1818_ngat), .B(G4658GAT_1744_ngat), .Y(G4896GAT_1847_gat) );
AND2XL U_g1817 (.A(G720GAT_228_ngat), .B(G4829GAT_1818_ngat), .Y(G4895GAT_1848_gat) );
AND2XL U_g1818 (.A(G4825GAT_1819_ngat), .B(G4654GAT_1745_ngat), .Y(G4891GAT_1849_gat) );
AND2XL U_g1819 (.A(G672GAT_244_ngat), .B(G4825GAT_1819_ngat), .Y(G4890GAT_1850_gat) );
AND2XL U_g1820 (.A(G4821GAT_1820_ngat), .B(G4650GAT_1746_ngat), .Y(G4886GAT_1851_gat) );
AND2XL U_g1821 (.A(G624GAT_260_ngat), .B(G4821GAT_1820_ngat), .Y(G4885GAT_1852_gat) );
AND2XL U_g1822 (.A(G4817GAT_1821_ngat), .B(G4646GAT_1747_ngat), .Y(G4881GAT_1853_gat) );
AND2XL U_g1823 (.A(G576GAT_276_ngat), .B(G4817GAT_1821_ngat), .Y(G4880GAT_1854_gat) );
AND2XL U_g1824 (.A(G4943GAT_1822_ngat), .B(G1302GAT_34_ngat), .Y(G5001GAT_1855_gat) );
AND2XL U_g1825 (.A(G4942GAT_1837_ngat), .B(G4941GAT_1823_ngat), .Y(G4998GAT_1856_gat) );
AND2XL U_g1826 (.A(G4937GAT_1839_ngat), .B(G4754GAT_1750_ngat), .Y(G4995GAT_1857_gat) );
AND2XL U_g1827 (.A(G4937GAT_1839_ngat), .B(G4872GAT_1799_ngat), .Y(G4993GAT_1858_gat) );
AND2XL U_g1828 (.A(G4933GAT_1826_ngat), .B(G4932GAT_1825_ngat), .Y(G4986GAT_1859_gat) );
AND2XL U_g1829 (.A(G4928GAT_1827_ngat), .B(G4863GAT_1803_ngat), .Y(G4984GAT_1860_gat) );
AND2XL U_g1830 (.A(G4860GAT_1804_ngat), .B(G4928GAT_1827_ngat), .Y(G4985GAT_1861_gat) );
AND2XL U_g1831 (.A(G4922GAT_1829_ngat), .B(G4925GAT_1828_ngat), .Y(G4980GAT_1862_gat) );
AND2XL U_g1832 (.A(G4921GAT_1843_ngat), .B(G4920GAT_1830_ngat), .Y(G4977GAT_1863_gat) );
AND2XL U_g1833 (.A(G4916GAT_1844_ngat), .B(G4733GAT_1757_ngat), .Y(G4974GAT_1864_gat) );
AND2XL U_g1834 (.A(G4916GAT_1844_ngat), .B(G4851GAT_1806_ngat), .Y(G4972GAT_1865_gat) );
AND2XL U_g1835 (.A(G4912GAT_1833_ngat), .B(G4911GAT_1832_ngat), .Y(G4965GAT_1866_gat) );
AND2XL U_g1836 (.A(G4907GAT_1834_ngat), .B(G4842GAT_1810_ngat), .Y(G4963GAT_1867_gat) );
AND2XL U_g1837 (.A(G4839GAT_1811_ngat), .B(G4907GAT_1834_ngat), .Y(G4964GAT_1868_gat) );
AND2XL U_g1838 (.A(G4901GAT_1845_ngat), .B(G4904GAT_1835_ngat), .Y(G4959GAT_1869_gat) );
AND2XL U_g1839 (.A(G4900GAT_1846_ngat), .B(G4899GAT_1836_ngat), .Y(G4956GAT_1870_gat) );
AND2XL U_g1840 (.A(G4895GAT_1848_ngat), .B(G4894GAT_1838_ngat), .Y(G4953GAT_1871_gat) );
AND2XL U_g1841 (.A(G1206GAT_66_ngat), .B(G4937GAT_1839_ngat), .Y(G4994GAT_1872_gat) );
AND2XL U_g1842 (.A(G4890GAT_1850_ngat), .B(G4889GAT_1840_ngat), .Y(G4950GAT_1873_gat) );
AND2XL U_g1843 (.A(G1158GAT_82_ngat), .B(G4934GAT_1824_ngat), .Y(G4989GAT_1874_gat) );
AND2XL U_g1844 (.A(G4885GAT_1852_ngat), .B(G4884GAT_1841_ngat), .Y(G4947GAT_1875_gat) );
AND2XL U_g1845 (.A(G4880GAT_1854_ngat), .B(G4879GAT_1842_ngat), .Y(G4946GAT_1876_gat) );
AND2XL U_g1846 (.A(G963GAT_147_ngat), .B(G4916GAT_1844_ngat), .Y(G4973GAT_1877_gat) );
AND2XL U_g1847 (.A(G915GAT_163_ngat), .B(G4913GAT_1831_ngat), .Y(G4968GAT_1878_gat) );
AND2XL U_g1848 (.A(G5001GAT_1855_ngat), .B(G1302GAT_34_ngat), .Y(G5063GAT_1879_gat) );
AND2XL U_g1849 (.A(G4943GAT_1822_ngat), .B(G5001GAT_1855_ngat), .Y(G5064GAT_1880_gat) );
AND2XL U_g1850 (.A(G4995GAT_1857_ngat), .B(G4998GAT_1856_ngat), .Y(G5059GAT_1881_gat) );
AND2XL U_g1851 (.A(G4994GAT_1872_ngat), .B(G4993GAT_1858_ngat), .Y(G5056GAT_1882_gat) );
AND2XL U_g1852 (.A(G4989GAT_1874_ngat), .B(G4808GAT_1779_ngat), .Y(G5053GAT_1883_gat) );
AND2XL U_g1853 (.A(G4989GAT_1874_ngat), .B(G4934GAT_1824_ngat), .Y(G5051GAT_1884_gat) );
AND2XL U_g1854 (.A(G4985GAT_1861_ngat), .B(G4984GAT_1860_ngat), .Y(G5044GAT_1885_gat) );
AND2XL U_g1855 (.A(G4980GAT_1862_ngat), .B(G4925GAT_1828_ngat), .Y(G5042GAT_1886_gat) );
AND2XL U_g1856 (.A(G4922GAT_1829_ngat), .B(G4980GAT_1862_ngat), .Y(G5043GAT_1887_gat) );
AND2XL U_g1857 (.A(G4974GAT_1864_ngat), .B(G4977GAT_1863_ngat), .Y(G5038GAT_1888_gat) );
AND2XL U_g1858 (.A(G4973GAT_1877_ngat), .B(G4972GAT_1865_ngat), .Y(G5035GAT_1889_gat) );
AND2XL U_g1859 (.A(G4968GAT_1878_ngat), .B(G4787GAT_1786_ngat), .Y(G5032GAT_1890_gat) );
AND2XL U_g1860 (.A(G4968GAT_1878_ngat), .B(G4913GAT_1831_ngat), .Y(G5030GAT_1891_gat) );
AND2XL U_g1861 (.A(G4964GAT_1868_ngat), .B(G4963GAT_1867_ngat), .Y(G5023GAT_1892_gat) );
AND2XL U_g1862 (.A(G4959GAT_1869_ngat), .B(G4904GAT_1835_ngat), .Y(G5021GAT_1893_gat) );
AND2XL U_g1863 (.A(G1158GAT_82_ngat), .B(G4989GAT_1874_ngat), .Y(G5052GAT_1894_gat) );
AND2XL U_g1864 (.A(G1110GAT_98_ngat), .B(G4986GAT_1859_ngat), .Y(G5047GAT_1895_gat) );
AND2XL U_g1865 (.A(G915GAT_163_ngat), .B(G4968GAT_1878_ngat), .Y(G5031GAT_1896_gat) );
AND2XL U_g1866 (.A(G867GAT_179_ngat), .B(G4965GAT_1866_ngat), .Y(G5026GAT_1897_gat) );
AND2XL U_g1867 (.A(G4901GAT_1845_ngat), .B(G4959GAT_1869_ngat), .Y(G5022GAT_1898_gat) );
AND2XL U_g1868 (.A(G4896GAT_1847_ngat), .B(G4956GAT_1870_ngat), .Y(G5017GAT_1899_gat) );
AND2XL U_g1869 (.A(G4891GAT_1849_ngat), .B(G4953GAT_1871_ngat), .Y(G5013GAT_1900_gat) );
AND2XL U_g1870 (.A(G4886GAT_1851_ngat), .B(G4950GAT_1873_ngat), .Y(G5009GAT_1901_gat) );
AND2XL U_g1871 (.A(G4881GAT_1853_ngat), .B(G4947GAT_1875_ngat), .Y(G5005GAT_1902_gat) );
AND2XL U_g1872 (.A(G5064GAT_1880_ngat), .B(G5063GAT_1879_ngat), .Y(G5115GAT_1903_gat) );
AND2XL U_g1873 (.A(G5059GAT_1881_ngat), .B(G4998GAT_1856_ngat), .Y(G5113GAT_1904_gat) );
AND2XL U_g1874 (.A(G4995GAT_1857_ngat), .B(G5059GAT_1881_ngat), .Y(G5114GAT_1905_gat) );
AND2XL U_g1875 (.A(G5053GAT_1883_ngat), .B(G5056GAT_1882_ngat), .Y(G5109GAT_1906_gat) );
AND2XL U_g1876 (.A(G5052GAT_1894_ngat), .B(G5051GAT_1884_ngat), .Y(G5106GAT_1907_gat) );
AND2XL U_g1877 (.A(G5047GAT_1895_ngat), .B(G4866GAT_1802_ngat), .Y(G5103GAT_1908_gat) );
AND2XL U_g1878 (.A(G5047GAT_1895_ngat), .B(G4986GAT_1859_ngat), .Y(G5101GAT_1909_gat) );
AND2XL U_g1879 (.A(G5043GAT_1887_ngat), .B(G5042GAT_1886_ngat), .Y(G5094GAT_1910_gat) );
AND2XL U_g1880 (.A(G5038GAT_1888_ngat), .B(G4977GAT_1863_ngat), .Y(G5092GAT_1911_gat) );
AND2XL U_g1881 (.A(G4974GAT_1864_ngat), .B(G5038GAT_1888_ngat), .Y(G5093GAT_1912_gat) );
AND2XL U_g1882 (.A(G5032GAT_1890_ngat), .B(G5035GAT_1889_ngat), .Y(G5088GAT_1913_gat) );
AND2XL U_g1883 (.A(G5031GAT_1896_ngat), .B(G5030GAT_1891_ngat), .Y(G5085GAT_1914_gat) );
AND2XL U_g1884 (.A(G5026GAT_1897_ngat), .B(G4845GAT_1809_ngat), .Y(G5082GAT_1915_gat) );
AND2XL U_g1885 (.A(G5026GAT_1897_ngat), .B(G4965GAT_1866_ngat), .Y(G5080GAT_1916_gat) );
AND2XL U_g1886 (.A(G5022GAT_1898_ngat), .B(G5021GAT_1893_ngat), .Y(G5073GAT_1917_gat) );
AND2XL U_g1887 (.A(G5017GAT_1899_ngat), .B(G4956GAT_1870_ngat), .Y(G5071GAT_1918_gat) );
AND2XL U_g1888 (.A(G5013GAT_1900_ngat), .B(G4953GAT_1871_ngat), .Y(G5069GAT_1919_gat) );
AND2XL U_g1889 (.A(G5009GAT_1901_ngat), .B(G4950GAT_1873_ngat), .Y(G5067GAT_1920_gat) );
AND2XL U_g1890 (.A(G5005GAT_1902_ngat), .B(G4947GAT_1875_ngat), .Y(G5065GAT_1921_gat) );
AND2XL U_g1891 (.A(G1110GAT_98_ngat), .B(G5047GAT_1895_ngat), .Y(G5102GAT_1922_gat) );
AND2XL U_g1892 (.A(G1062GAT_114_ngat), .B(G5044GAT_1885_ngat), .Y(G5097GAT_1923_gat) );
AND2XL U_g1893 (.A(G867GAT_179_ngat), .B(G5026GAT_1897_ngat), .Y(G5081GAT_1924_gat) );
AND2XL U_g1894 (.A(G819GAT_195_ngat), .B(G5023GAT_1892_ngat), .Y(G5076GAT_1925_gat) );
AND2XL U_g1895 (.A(G4896GAT_1847_ngat), .B(G5017GAT_1899_ngat), .Y(G5072GAT_1926_gat) );
AND2XL U_g1896 (.A(G4891GAT_1849_ngat), .B(G5013GAT_1900_ngat), .Y(G5070GAT_1927_gat) );
AND2XL U_g1897 (.A(G4886GAT_1851_ngat), .B(G5009GAT_1901_ngat), .Y(G5068GAT_1928_gat) );
AND2XL U_g1898 (.A(G4881GAT_1853_ngat), .B(G5005GAT_1902_ngat), .Y(G5066GAT_1929_gat) );
AND2XL U_g1899 (.A(G5114GAT_1905_ngat), .B(G5113GAT_1904_ngat), .Y(G5169GAT_1930_gat) );
AND2XL U_g1900 (.A(G5109GAT_1906_ngat), .B(G5056GAT_1882_ngat), .Y(G5167GAT_1931_gat) );
AND2XL U_g1901 (.A(G5053GAT_1883_ngat), .B(G5109GAT_1906_ngat), .Y(G5168GAT_1932_gat) );
AND2XL U_g1902 (.A(G5103GAT_1908_ngat), .B(G5106GAT_1907_ngat), .Y(G5163GAT_1933_gat) );
AND2XL U_g1903 (.A(G5102GAT_1922_ngat), .B(G5101GAT_1909_ngat), .Y(G5160GAT_1934_gat) );
AND2XL U_g1904 (.A(G5097GAT_1923_ngat), .B(G4928GAT_1827_ngat), .Y(G5157GAT_1935_gat) );
AND2XL U_g1905 (.A(G5097GAT_1923_ngat), .B(G5044GAT_1885_ngat), .Y(G5155GAT_1936_gat) );
AND2XL U_g1906 (.A(G5093GAT_1912_ngat), .B(G5092GAT_1911_ngat), .Y(G5148GAT_1937_gat) );
AND2XL U_g1907 (.A(G5088GAT_1913_ngat), .B(G5035GAT_1889_ngat), .Y(G5146GAT_1938_gat) );
AND2XL U_g1908 (.A(G5032GAT_1890_ngat), .B(G5088GAT_1913_ngat), .Y(G5147GAT_1939_gat) );
AND2XL U_g1909 (.A(G5082GAT_1915_ngat), .B(G5085GAT_1914_ngat), .Y(G5142GAT_1940_gat) );
AND2XL U_g1910 (.A(G5081GAT_1924_ngat), .B(G5080GAT_1916_ngat), .Y(G5139GAT_1941_gat) );
AND2XL U_g1911 (.A(G5076GAT_1925_ngat), .B(G4907GAT_1834_ngat), .Y(G5136GAT_1942_gat) );
AND2XL U_g1912 (.A(G5076GAT_1925_ngat), .B(G5023GAT_1892_ngat), .Y(G5134GAT_1943_gat) );
AND2XL U_g1913 (.A(G5072GAT_1926_ngat), .B(G5071GAT_1918_ngat), .Y(G5127GAT_1944_gat) );
AND2XL U_g1914 (.A(G1257GAT_49_ngat), .B(G5115GAT_1903_ngat), .Y(G5172GAT_1945_gat) );
AND2XL U_g1915 (.A(G5070GAT_1927_ngat), .B(G5069GAT_1919_ngat), .Y(G5124GAT_1946_gat) );
AND2XL U_g1916 (.A(G5068GAT_1928_ngat), .B(G5067GAT_1920_ngat), .Y(G5121GAT_1947_gat) );
AND2XL U_g1917 (.A(G5066GAT_1929_ngat), .B(G5065GAT_1921_ngat), .Y(G5118GAT_1948_gat) );
AND2XL U_g1918 (.A(G1062GAT_114_ngat), .B(G5097GAT_1923_ngat), .Y(G5156GAT_1949_gat) );
AND2XL U_g1919 (.A(G1014GAT_130_ngat), .B(G5094GAT_1910_ngat), .Y(G5151GAT_1950_gat) );
AND2XL U_g1920 (.A(G819GAT_195_ngat), .B(G5076GAT_1925_ngat), .Y(G5135GAT_1951_gat) );
AND2XL U_g1921 (.A(G771GAT_211_ngat), .B(G5073GAT_1917_ngat), .Y(G5130GAT_1952_gat) );
AND2XL U_g1922 (.A(G5172GAT_1945_ngat), .B(G5001GAT_1855_ngat), .Y(G5236GAT_1953_gat) );
AND2XL U_g1923 (.A(G5172GAT_1945_ngat), .B(G5115GAT_1903_ngat), .Y(G5234GAT_1954_gat) );
AND2XL U_g1924 (.A(G5168GAT_1932_ngat), .B(G5167GAT_1931_ngat), .Y(G5227GAT_1955_gat) );
AND2XL U_g1925 (.A(G5163GAT_1933_ngat), .B(G5106GAT_1907_ngat), .Y(G5225GAT_1956_gat) );
AND2XL U_g1926 (.A(G5103GAT_1908_ngat), .B(G5163GAT_1933_ngat), .Y(G5226GAT_1957_gat) );
AND2XL U_g1927 (.A(G5157GAT_1935_ngat), .B(G5160GAT_1934_ngat), .Y(G5221GAT_1958_gat) );
AND2XL U_g1928 (.A(G5156GAT_1949_ngat), .B(G5155GAT_1936_ngat), .Y(G5218GAT_1959_gat) );
AND2XL U_g1929 (.A(G5151GAT_1950_ngat), .B(G4980GAT_1862_ngat), .Y(G5215GAT_1960_gat) );
AND2XL U_g1930 (.A(G5151GAT_1950_ngat), .B(G5094GAT_1910_ngat), .Y(G5213GAT_1961_gat) );
AND2XL U_g1931 (.A(G5147GAT_1939_ngat), .B(G5146GAT_1938_ngat), .Y(G5206GAT_1962_gat) );
AND2XL U_g1932 (.A(G5142GAT_1940_ngat), .B(G5085GAT_1914_ngat), .Y(G5204GAT_1963_gat) );
AND2XL U_g1933 (.A(G5082GAT_1915_ngat), .B(G5142GAT_1940_ngat), .Y(G5205GAT_1964_gat) );
AND2XL U_g1934 (.A(G5136GAT_1942_ngat), .B(G5139GAT_1941_ngat), .Y(G5200GAT_1965_gat) );
AND2XL U_g1935 (.A(G5135GAT_1951_ngat), .B(G5134GAT_1943_ngat), .Y(G5197GAT_1966_gat) );
AND2XL U_g1936 (.A(G5130GAT_1952_ngat), .B(G4959GAT_1869_ngat), .Y(G5194GAT_1967_gat) );
AND2XL U_g1937 (.A(G5130GAT_1952_ngat), .B(G5073GAT_1917_ngat), .Y(G5192GAT_1968_gat) );
AND2XL U_g1938 (.A(G1257GAT_49_ngat), .B(G5172GAT_1945_ngat), .Y(G5235GAT_1969_gat) );
AND2XL U_g1939 (.A(G1209GAT_65_ngat), .B(G5169GAT_1930_ngat), .Y(G5230GAT_1970_gat) );
AND2XL U_g1940 (.A(G1014GAT_130_ngat), .B(G5151GAT_1950_ngat), .Y(G5214GAT_1971_gat) );
AND2XL U_g1941 (.A(G966GAT_146_ngat), .B(G5148GAT_1937_ngat), .Y(G5209GAT_1972_gat) );
AND2XL U_g1942 (.A(G771GAT_211_ngat), .B(G5130GAT_1952_ngat), .Y(G5193GAT_1973_gat) );
AND2XL U_g1943 (.A(G723GAT_227_ngat), .B(G5127GAT_1944_ngat), .Y(G5188GAT_1974_gat) );
AND2XL U_g1944 (.A(G675GAT_243_ngat), .B(G5124GAT_1946_ngat), .Y(G5184GAT_1975_gat) );
AND2XL U_g1945 (.A(G627GAT_259_ngat), .B(G5121GAT_1947_ngat), .Y(G5180GAT_1976_gat) );
AND2XL U_g1946 (.A(G579GAT_275_ngat), .B(G5118GAT_1948_ngat), .Y(G5176GAT_1977_gat) );
AND2XL U_g1947 (.A(G5236GAT_1953_ngat), .B(G1305GAT_33_ngat), .Y(G5304GAT_1978_gat) );
AND2XL U_g1948 (.A(G5235GAT_1969_ngat), .B(G5234GAT_1954_ngat), .Y(G5301GAT_1979_gat) );
AND2XL U_g1949 (.A(G5230GAT_1970_ngat), .B(G5059GAT_1881_ngat), .Y(G5298GAT_1980_gat) );
AND2XL U_g1950 (.A(G5230GAT_1970_ngat), .B(G5169GAT_1930_ngat), .Y(G5296GAT_1981_gat) );
AND2XL U_g1951 (.A(G5226GAT_1957_ngat), .B(G5225GAT_1956_ngat), .Y(G5289GAT_1982_gat) );
AND2XL U_g1952 (.A(G5221GAT_1958_ngat), .B(G5160GAT_1934_ngat), .Y(G5287GAT_1983_gat) );
AND2XL U_g1953 (.A(G5157GAT_1935_ngat), .B(G5221GAT_1958_ngat), .Y(G5288GAT_1984_gat) );
AND2XL U_g1954 (.A(G5215GAT_1960_ngat), .B(G5218GAT_1959_ngat), .Y(G5283GAT_1985_gat) );
AND2XL U_g1955 (.A(G5214GAT_1971_ngat), .B(G5213GAT_1961_ngat), .Y(G5280GAT_1986_gat) );
AND2XL U_g1956 (.A(G5209GAT_1972_ngat), .B(G5038GAT_1888_ngat), .Y(G5277GAT_1987_gat) );
AND2XL U_g1957 (.A(G5209GAT_1972_ngat), .B(G5148GAT_1937_ngat), .Y(G5275GAT_1988_gat) );
AND2XL U_g1958 (.A(G5205GAT_1964_ngat), .B(G5204GAT_1963_ngat), .Y(G5268GAT_1989_gat) );
AND2XL U_g1959 (.A(G5200GAT_1965_ngat), .B(G5139GAT_1941_ngat), .Y(G5266GAT_1990_gat) );
AND2XL U_g1960 (.A(G5136GAT_1942_ngat), .B(G5200GAT_1965_ngat), .Y(G5267GAT_1991_gat) );
AND2XL U_g1961 (.A(G5194GAT_1967_ngat), .B(G5197GAT_1966_ngat), .Y(G5262GAT_1992_gat) );
AND2XL U_g1962 (.A(G5193GAT_1973_ngat), .B(G5192GAT_1968_ngat), .Y(G5259GAT_1993_gat) );
AND2XL U_g1963 (.A(G5188GAT_1974_ngat), .B(G5127GAT_1944_ngat), .Y(G5254GAT_1994_gat) );
AND2XL U_g1964 (.A(G5184GAT_1975_ngat), .B(G5124GAT_1946_ngat), .Y(G5249GAT_1995_gat) );
AND2XL U_g1965 (.A(G1209GAT_65_ngat), .B(G5230GAT_1970_ngat), .Y(G5297GAT_1996_gat) );
AND2XL U_g1966 (.A(G5180GAT_1976_ngat), .B(G5121GAT_1947_ngat), .Y(G5244GAT_1997_gat) );
AND2XL U_g1967 (.A(G1161GAT_81_ngat), .B(G5227GAT_1955_ngat), .Y(G5292GAT_1998_gat) );
AND2XL U_g1968 (.A(G5176GAT_1977_ngat), .B(G5118GAT_1948_ngat), .Y(G5239GAT_1999_gat) );
AND2XL U_g1969 (.A(G966GAT_146_ngat), .B(G5209GAT_1972_ngat), .Y(G5276GAT_2000_gat) );
AND2XL U_g1970 (.A(G918GAT_162_ngat), .B(G5206GAT_1962_ngat), .Y(G5271GAT_2001_gat) );
AND2XL U_g1971 (.A(G5188GAT_1974_ngat), .B(G5017GAT_1899_ngat), .Y(G5256GAT_2002_gat) );
AND2XL U_g1972 (.A(G723GAT_227_ngat), .B(G5188GAT_1974_ngat), .Y(G5255GAT_2003_gat) );
AND2XL U_g1973 (.A(G5184GAT_1975_ngat), .B(G5013GAT_1900_ngat), .Y(G5251GAT_2004_gat) );
AND2XL U_g1974 (.A(G675GAT_243_ngat), .B(G5184GAT_1975_ngat), .Y(G5250GAT_2005_gat) );
AND2XL U_g1975 (.A(G5180GAT_1976_ngat), .B(G5009GAT_1901_ngat), .Y(G5246GAT_2006_gat) );
AND2XL U_g1976 (.A(G627GAT_259_ngat), .B(G5180GAT_1976_ngat), .Y(G5245GAT_2007_gat) );
AND2XL U_g1977 (.A(G5176GAT_1977_ngat), .B(G5005GAT_1902_ngat), .Y(G5241GAT_2008_gat) );
AND2XL U_g1978 (.A(G579GAT_275_ngat), .B(G5176GAT_1977_ngat), .Y(G5240GAT_2009_gat) );
AND2XL U_g1979 (.A(G5304GAT_1978_ngat), .B(G1305GAT_33_ngat), .Y(G5364GAT_2010_gat) );
AND2XL U_g1980 (.A(G5236GAT_1953_ngat), .B(G5304GAT_1978_ngat), .Y(G5365GAT_2011_gat) );
AND2XL U_g1981 (.A(G5298GAT_1980_ngat), .B(G5301GAT_1979_ngat), .Y(G5360GAT_2012_gat) );
AND2XL U_g1982 (.A(G5297GAT_1996_ngat), .B(G5296GAT_1981_ngat), .Y(G5357GAT_2013_gat) );
AND2XL U_g1983 (.A(G5292GAT_1998_ngat), .B(G5109GAT_1906_ngat), .Y(G5354GAT_2014_gat) );
AND2XL U_g1984 (.A(G5292GAT_1998_ngat), .B(G5227GAT_1955_ngat), .Y(G5352GAT_2015_gat) );
AND2XL U_g1985 (.A(G5288GAT_1984_ngat), .B(G5287GAT_1983_ngat), .Y(G5345GAT_2016_gat) );
AND2XL U_g1986 (.A(G5283GAT_1985_ngat), .B(G5218GAT_1959_ngat), .Y(G5343GAT_2017_gat) );
AND2XL U_g1987 (.A(G5215GAT_1960_ngat), .B(G5283GAT_1985_ngat), .Y(G5344GAT_2018_gat) );
AND2XL U_g1988 (.A(G5277GAT_1987_ngat), .B(G5280GAT_1986_ngat), .Y(G5339GAT_2019_gat) );
AND2XL U_g1989 (.A(G5276GAT_2000_ngat), .B(G5275GAT_1988_ngat), .Y(G5336GAT_2020_gat) );
AND2XL U_g1990 (.A(G5271GAT_2001_ngat), .B(G5088GAT_1913_ngat), .Y(G5333GAT_2021_gat) );
AND2XL U_g1991 (.A(G5271GAT_2001_ngat), .B(G5206GAT_1962_ngat), .Y(G5331GAT_2022_gat) );
AND2XL U_g1992 (.A(G5267GAT_1991_ngat), .B(G5266GAT_1990_ngat), .Y(G5324GAT_2023_gat) );
AND2XL U_g1993 (.A(G5262GAT_1992_ngat), .B(G5197GAT_1966_ngat), .Y(G5322GAT_2024_gat) );
AND2XL U_g1994 (.A(G5194GAT_1967_ngat), .B(G5262GAT_1992_ngat), .Y(G5323GAT_2025_gat) );
AND2XL U_g1995 (.A(G5256GAT_2002_ngat), .B(G5259GAT_1993_ngat), .Y(G5318GAT_2026_gat) );
AND2XL U_g1996 (.A(G5255GAT_2003_ngat), .B(G5254GAT_1994_ngat), .Y(G5315GAT_2027_gat) );
AND2XL U_g1997 (.A(G5250GAT_2005_ngat), .B(G5249GAT_1995_ngat), .Y(G5312GAT_2028_gat) );
AND2XL U_g1998 (.A(G5245GAT_2007_ngat), .B(G5244GAT_1997_ngat), .Y(G5309GAT_2029_gat) );
AND2XL U_g1999 (.A(G1161GAT_81_ngat), .B(G5292GAT_1998_ngat), .Y(G5353GAT_2030_gat) );
AND2XL U_g2000 (.A(G5240GAT_2009_ngat), .B(G5239GAT_1999_ngat), .Y(G5308GAT_2031_gat) );
AND2XL U_g2001 (.A(G1113GAT_97_ngat), .B(G5289GAT_1982_ngat), .Y(G5348GAT_2032_gat) );
AND2XL U_g2002 (.A(G918GAT_162_ngat), .B(G5271GAT_2001_ngat), .Y(G5332GAT_2033_gat) );
AND2XL U_g2003 (.A(G870GAT_178_ngat), .B(G5268GAT_1989_ngat), .Y(G5327GAT_2034_gat) );
AND2XL U_g2004 (.A(G5365GAT_2011_ngat), .B(G5364GAT_2010_ngat), .Y(G5422GAT_2035_gat) );
AND2XL U_g2005 (.A(G5360GAT_2012_ngat), .B(G5301GAT_1979_ngat), .Y(G5420GAT_2036_gat) );
AND2XL U_g2006 (.A(G5298GAT_1980_ngat), .B(G5360GAT_2012_ngat), .Y(G5421GAT_2037_gat) );
AND2XL U_g2007 (.A(G5354GAT_2014_ngat), .B(G5357GAT_2013_ngat), .Y(G5416GAT_2038_gat) );
AND2XL U_g2008 (.A(G5353GAT_2030_ngat), .B(G5352GAT_2015_ngat), .Y(G5413GAT_2039_gat) );
AND2XL U_g2009 (.A(G5348GAT_2032_ngat), .B(G5163GAT_1933_ngat), .Y(G5410GAT_2040_gat) );
AND2XL U_g2010 (.A(G5348GAT_2032_ngat), .B(G5289GAT_1982_ngat), .Y(G5408GAT_2041_gat) );
AND2XL U_g2011 (.A(G5344GAT_2018_ngat), .B(G5343GAT_2017_ngat), .Y(G5401GAT_2042_gat) );
AND2XL U_g2012 (.A(G5339GAT_2019_ngat), .B(G5280GAT_1986_ngat), .Y(G5399GAT_2043_gat) );
AND2XL U_g2013 (.A(G5277GAT_1987_ngat), .B(G5339GAT_2019_ngat), .Y(G5400GAT_2044_gat) );
AND2XL U_g2014 (.A(G5333GAT_2021_ngat), .B(G5336GAT_2020_ngat), .Y(G5395GAT_2045_gat) );
AND2XL U_g2015 (.A(G5332GAT_2033_ngat), .B(G5331GAT_2022_ngat), .Y(G5392GAT_2046_gat) );
AND2XL U_g2016 (.A(G5327GAT_2034_ngat), .B(G5142GAT_1940_ngat), .Y(G5389GAT_2047_gat) );
AND2XL U_g2017 (.A(G5327GAT_2034_ngat), .B(G5268GAT_1989_ngat), .Y(G5387GAT_2048_gat) );
AND2XL U_g2018 (.A(G5323GAT_2025_ngat), .B(G5322GAT_2024_ngat), .Y(G5380GAT_2049_gat) );
AND2XL U_g2019 (.A(G5318GAT_2026_ngat), .B(G5259GAT_1993_ngat), .Y(G5378GAT_2050_gat) );
AND2XL U_g2020 (.A(G1113GAT_97_ngat), .B(G5348GAT_2032_ngat), .Y(G5409GAT_2051_gat) );
AND2XL U_g2021 (.A(G1065GAT_113_ngat), .B(G5345GAT_2016_ngat), .Y(G5404GAT_2052_gat) );
AND2XL U_g2022 (.A(G870GAT_178_ngat), .B(G5327GAT_2034_ngat), .Y(G5388GAT_2053_gat) );
AND2XL U_g2023 (.A(G822GAT_194_ngat), .B(G5324GAT_2023_ngat), .Y(G5383GAT_2054_gat) );
AND2XL U_g2024 (.A(G5256GAT_2002_ngat), .B(G5318GAT_2026_ngat), .Y(G5379GAT_2055_gat) );
AND2XL U_g2025 (.A(G5251GAT_2004_ngat), .B(G5315GAT_2027_ngat), .Y(G5374GAT_2056_gat) );
AND2XL U_g2026 (.A(G5246GAT_2006_ngat), .B(G5312GAT_2028_ngat), .Y(G5370GAT_2057_gat) );
AND2XL U_g2027 (.A(G5241GAT_2008_ngat), .B(G5309GAT_2029_ngat), .Y(G5366GAT_2058_gat) );
AND2XL U_g2028 (.A(G5421GAT_2037_ngat), .B(G5420GAT_2036_ngat), .Y(G5473GAT_2059_gat) );
AND2XL U_g2029 (.A(G5416GAT_2038_ngat), .B(G5357GAT_2013_ngat), .Y(G5471GAT_2060_gat) );
AND2XL U_g2030 (.A(G5354GAT_2014_ngat), .B(G5416GAT_2038_ngat), .Y(G5472GAT_2061_gat) );
AND2XL U_g2031 (.A(G5410GAT_2040_ngat), .B(G5413GAT_2039_ngat), .Y(G5467GAT_2062_gat) );
AND2XL U_g2032 (.A(G5409GAT_2051_ngat), .B(G5408GAT_2041_ngat), .Y(G5464GAT_2063_gat) );
AND2XL U_g2033 (.A(G5404GAT_2052_ngat), .B(G5221GAT_1958_ngat), .Y(G5461GAT_2064_gat) );
AND2XL U_g2034 (.A(G5404GAT_2052_ngat), .B(G5345GAT_2016_ngat), .Y(G5459GAT_2065_gat) );
AND2XL U_g2035 (.A(G5400GAT_2044_ngat), .B(G5399GAT_2043_ngat), .Y(G5452GAT_2066_gat) );
AND2XL U_g2036 (.A(G5395GAT_2045_ngat), .B(G5336GAT_2020_ngat), .Y(G5450GAT_2067_gat) );
AND2XL U_g2037 (.A(G5333GAT_2021_ngat), .B(G5395GAT_2045_ngat), .Y(G5451GAT_2068_gat) );
AND2XL U_g2038 (.A(G5389GAT_2047_ngat), .B(G5392GAT_2046_ngat), .Y(G5446GAT_2069_gat) );
AND2XL U_g2039 (.A(G5388GAT_2053_ngat), .B(G5387GAT_2048_ngat), .Y(G5443GAT_2070_gat) );
AND2XL U_g2040 (.A(G5383GAT_2054_ngat), .B(G5200GAT_1965_ngat), .Y(G5440GAT_2071_gat) );
AND2XL U_g2041 (.A(G5383GAT_2054_ngat), .B(G5324GAT_2023_ngat), .Y(G5438GAT_2072_gat) );
AND2XL U_g2042 (.A(G5379GAT_2055_ngat), .B(G5378GAT_2050_ngat), .Y(G5431GAT_2073_gat) );
AND2XL U_g2043 (.A(G5374GAT_2056_ngat), .B(G5315GAT_2027_ngat), .Y(G5429GAT_2074_gat) );
AND2XL U_g2044 (.A(G1260GAT_48_ngat), .B(G5422GAT_2035_ngat), .Y(G5476GAT_2075_gat) );
AND2XL U_g2045 (.A(G5370GAT_2057_ngat), .B(G5312GAT_2028_ngat), .Y(G5427GAT_2076_gat) );
AND2XL U_g2046 (.A(G5366GAT_2058_ngat), .B(G5309GAT_2029_ngat), .Y(G5425GAT_2077_gat) );
AND2XL U_g2047 (.A(G1065GAT_113_ngat), .B(G5404GAT_2052_ngat), .Y(G5460GAT_2078_gat) );
AND2XL U_g2048 (.A(G1017GAT_129_ngat), .B(G5401GAT_2042_ngat), .Y(G5455GAT_2079_gat) );
AND2XL U_g2049 (.A(G822GAT_194_ngat), .B(G5383GAT_2054_ngat), .Y(G5439GAT_2080_gat) );
AND2XL U_g2050 (.A(G774GAT_210_ngat), .B(G5380GAT_2049_ngat), .Y(G5434GAT_2081_gat) );
AND2XL U_g2051 (.A(G5251GAT_2004_ngat), .B(G5374GAT_2056_ngat), .Y(G5430GAT_2082_gat) );
AND2XL U_g2052 (.A(G5246GAT_2006_ngat), .B(G5370GAT_2057_ngat), .Y(G5428GAT_2083_gat) );
AND2XL U_g2053 (.A(G5241GAT_2008_ngat), .B(G5366GAT_2058_ngat), .Y(G5426GAT_2084_gat) );
AND2XL U_g2054 (.A(G5476GAT_2075_ngat), .B(G5304GAT_1978_ngat), .Y(G5537GAT_2085_gat) );
AND2XL U_g2055 (.A(G5476GAT_2075_ngat), .B(G5422GAT_2035_ngat), .Y(G5535GAT_2086_gat) );
AND2XL U_g2056 (.A(G5472GAT_2061_ngat), .B(G5471GAT_2060_ngat), .Y(G5528GAT_2087_gat) );
AND2XL U_g2057 (.A(G5467GAT_2062_ngat), .B(G5413GAT_2039_ngat), .Y(G5526GAT_2088_gat) );
AND2XL U_g2058 (.A(G5410GAT_2040_ngat), .B(G5467GAT_2062_ngat), .Y(G5527GAT_2089_gat) );
AND2XL U_g2059 (.A(G5461GAT_2064_ngat), .B(G5464GAT_2063_ngat), .Y(G5522GAT_2090_gat) );
AND2XL U_g2060 (.A(G5460GAT_2078_ngat), .B(G5459GAT_2065_ngat), .Y(G5519GAT_2091_gat) );
AND2XL U_g2061 (.A(G5455GAT_2079_ngat), .B(G5283GAT_1985_ngat), .Y(G5516GAT_2092_gat) );
AND2XL U_g2062 (.A(G5455GAT_2079_ngat), .B(G5401GAT_2042_ngat), .Y(G5514GAT_2093_gat) );
AND2XL U_g2063 (.A(G5451GAT_2068_ngat), .B(G5450GAT_2067_ngat), .Y(G5507GAT_2094_gat) );
AND2XL U_g2064 (.A(G5446GAT_2069_ngat), .B(G5392GAT_2046_ngat), .Y(G5505GAT_2095_gat) );
AND2XL U_g2065 (.A(G5389GAT_2047_ngat), .B(G5446GAT_2069_ngat), .Y(G5506GAT_2096_gat) );
AND2XL U_g2066 (.A(G5440GAT_2071_ngat), .B(G5443GAT_2070_ngat), .Y(G5501GAT_2097_gat) );
AND2XL U_g2067 (.A(G5439GAT_2080_ngat), .B(G5438GAT_2072_ngat), .Y(G5498GAT_2098_gat) );
AND2XL U_g2068 (.A(G5434GAT_2081_ngat), .B(G5262GAT_1992_ngat), .Y(G5495GAT_2099_gat) );
AND2XL U_g2069 (.A(G5434GAT_2081_ngat), .B(G5380GAT_2049_ngat), .Y(G5493GAT_2100_gat) );
AND2XL U_g2070 (.A(G5430GAT_2082_ngat), .B(G5429GAT_2074_ngat), .Y(G5486GAT_2101_gat) );
AND2XL U_g2071 (.A(G1260GAT_48_ngat), .B(G5476GAT_2075_ngat), .Y(G5536GAT_2102_gat) );
AND2XL U_g2072 (.A(G5428GAT_2083_ngat), .B(G5427GAT_2076_ngat), .Y(G5483GAT_2103_gat) );
AND2XL U_g2073 (.A(G1212GAT_64_ngat), .B(G5473GAT_2059_ngat), .Y(G5531GAT_2104_gat) );
AND2XL U_g2074 (.A(G5426GAT_2084_ngat), .B(G5425GAT_2077_ngat), .Y(G5480GAT_2105_gat) );
AND2XL U_g2075 (.A(G1017GAT_129_ngat), .B(G5455GAT_2079_ngat), .Y(G5515GAT_2106_gat) );
AND2XL U_g2076 (.A(G969GAT_145_ngat), .B(G5452GAT_2066_ngat), .Y(G5510GAT_2107_gat) );
AND2XL U_g2077 (.A(G774GAT_210_ngat), .B(G5434GAT_2081_ngat), .Y(G5494GAT_2108_gat) );
AND2XL U_g2078 (.A(G726GAT_226_ngat), .B(G5431GAT_2073_ngat), .Y(G5489GAT_2109_gat) );
AND2XL U_g2079 (.A(G5537GAT_2085_ngat), .B(G1308GAT_32_ngat), .Y(G5602GAT_2110_gat) );
AND2XL U_g2080 (.A(G5536GAT_2102_ngat), .B(G5535GAT_2086_ngat), .Y(G5599GAT_2111_gat) );
AND2XL U_g2081 (.A(G5531GAT_2104_ngat), .B(G5360GAT_2012_ngat), .Y(G5596GAT_2112_gat) );
AND2XL U_g2082 (.A(G5531GAT_2104_ngat), .B(G5473GAT_2059_ngat), .Y(G5594GAT_2113_gat) );
AND2XL U_g2083 (.A(G5527GAT_2089_ngat), .B(G5526GAT_2088_ngat), .Y(G5587GAT_2114_gat) );
AND2XL U_g2084 (.A(G5522GAT_2090_ngat), .B(G5464GAT_2063_ngat), .Y(G5585GAT_2115_gat) );
AND2XL U_g2085 (.A(G5461GAT_2064_ngat), .B(G5522GAT_2090_ngat), .Y(G5586GAT_2116_gat) );
AND2XL U_g2086 (.A(G5516GAT_2092_ngat), .B(G5519GAT_2091_ngat), .Y(G5581GAT_2117_gat) );
AND2XL U_g2087 (.A(G5515GAT_2106_ngat), .B(G5514GAT_2093_ngat), .Y(G5578GAT_2118_gat) );
AND2XL U_g2088 (.A(G5510GAT_2107_ngat), .B(G5339GAT_2019_ngat), .Y(G5575GAT_2119_gat) );
AND2XL U_g2089 (.A(G5510GAT_2107_ngat), .B(G5452GAT_2066_ngat), .Y(G5573GAT_2120_gat) );
AND2XL U_g2090 (.A(G5506GAT_2096_ngat), .B(G5505GAT_2095_ngat), .Y(G5566GAT_2121_gat) );
AND2XL U_g2091 (.A(G5501GAT_2097_ngat), .B(G5443GAT_2070_ngat), .Y(G5564GAT_2122_gat) );
AND2XL U_g2092 (.A(G5440GAT_2071_ngat), .B(G5501GAT_2097_ngat), .Y(G5565GAT_2123_gat) );
AND2XL U_g2093 (.A(G5495GAT_2099_ngat), .B(G5498GAT_2098_ngat), .Y(G5560GAT_2124_gat) );
AND2XL U_g2094 (.A(G5494GAT_2108_ngat), .B(G5493GAT_2100_ngat), .Y(G5557GAT_2125_gat) );
AND2XL U_g2095 (.A(G5489GAT_2109_ngat), .B(G5318GAT_2026_ngat), .Y(G5554GAT_2126_gat) );
AND2XL U_g2096 (.A(G5489GAT_2109_ngat), .B(G5431GAT_2073_ngat), .Y(G5552GAT_2127_gat) );
AND2XL U_g2097 (.A(G1212GAT_64_ngat), .B(G5531GAT_2104_ngat), .Y(G5595GAT_2128_gat) );
AND2XL U_g2098 (.A(G1164GAT_80_ngat), .B(G5528GAT_2087_ngat), .Y(G5590GAT_2129_gat) );
AND2XL U_g2099 (.A(G969GAT_145_ngat), .B(G5510GAT_2107_ngat), .Y(G5574GAT_2130_gat) );
AND2XL U_g2100 (.A(G921GAT_161_ngat), .B(G5507GAT_2094_ngat), .Y(G5569GAT_2131_gat) );
AND2XL U_g2101 (.A(G726GAT_226_ngat), .B(G5489GAT_2109_ngat), .Y(G5553GAT_2132_gat) );
AND2XL U_g2102 (.A(G678GAT_242_ngat), .B(G5486GAT_2101_ngat), .Y(G5548GAT_2133_gat) );
AND2XL U_g2103 (.A(G630GAT_258_ngat), .B(G5483GAT_2103_ngat), .Y(G5544GAT_2134_gat) );
AND2XL U_g2104 (.A(G582GAT_274_ngat), .B(G5480GAT_2105_ngat), .Y(G5540GAT_2135_gat) );
AND2XL U_g2105 (.A(G5602GAT_2110_ngat), .B(G1308GAT_32_ngat), .Y(G5670GAT_2136_gat) );
AND2XL U_g2106 (.A(G5537GAT_2085_ngat), .B(G5602GAT_2110_ngat), .Y(G5671GAT_2137_gat) );
AND2XL U_g2107 (.A(G5596GAT_2112_ngat), .B(G5599GAT_2111_ngat), .Y(G5666GAT_2138_gat) );
AND2XL U_g2108 (.A(G5595GAT_2128_ngat), .B(G5594GAT_2113_ngat), .Y(G5663GAT_2139_gat) );
AND2XL U_g2109 (.A(G5590GAT_2129_ngat), .B(G5416GAT_2038_ngat), .Y(G5660GAT_2140_gat) );
AND2XL U_g2110 (.A(G5590GAT_2129_ngat), .B(G5528GAT_2087_ngat), .Y(G5658GAT_2141_gat) );
AND2XL U_g2111 (.A(G5586GAT_2116_ngat), .B(G5585GAT_2115_ngat), .Y(G5651GAT_2142_gat) );
AND2XL U_g2112 (.A(G5581GAT_2117_ngat), .B(G5519GAT_2091_ngat), .Y(G5649GAT_2143_gat) );
AND2XL U_g2113 (.A(G5516GAT_2092_ngat), .B(G5581GAT_2117_ngat), .Y(G5650GAT_2144_gat) );
AND2XL U_g2114 (.A(G5575GAT_2119_ngat), .B(G5578GAT_2118_ngat), .Y(G5645GAT_2145_gat) );
AND2XL U_g2115 (.A(G5574GAT_2130_ngat), .B(G5573GAT_2120_ngat), .Y(G5642GAT_2146_gat) );
AND2XL U_g2116 (.A(G5569GAT_2131_ngat), .B(G5395GAT_2045_ngat), .Y(G5639GAT_2147_gat) );
AND2XL U_g2117 (.A(G5569GAT_2131_ngat), .B(G5507GAT_2094_ngat), .Y(G5637GAT_2148_gat) );
AND2XL U_g2118 (.A(G5565GAT_2123_ngat), .B(G5564GAT_2122_ngat), .Y(G5630GAT_2149_gat) );
AND2XL U_g2119 (.A(G5560GAT_2124_ngat), .B(G5498GAT_2098_ngat), .Y(G5628GAT_2150_gat) );
AND2XL U_g2120 (.A(G5495GAT_2099_ngat), .B(G5560GAT_2124_ngat), .Y(G5629GAT_2151_gat) );
AND2XL U_g2121 (.A(G5554GAT_2126_ngat), .B(G5557GAT_2125_ngat), .Y(G5624GAT_2152_gat) );
AND2XL U_g2122 (.A(G5553GAT_2132_ngat), .B(G5552GAT_2127_ngat), .Y(G5621GAT_2153_gat) );
AND2XL U_g2123 (.A(G5548GAT_2133_ngat), .B(G5486GAT_2101_ngat), .Y(G5616GAT_2154_gat) );
AND2XL U_g2124 (.A(G5544GAT_2134_ngat), .B(G5483GAT_2103_ngat), .Y(G5611GAT_2155_gat) );
AND2XL U_g2125 (.A(G5540GAT_2135_ngat), .B(G5480GAT_2105_ngat), .Y(G5606GAT_2156_gat) );
AND2XL U_g2126 (.A(G1164GAT_80_ngat), .B(G5590GAT_2129_ngat), .Y(G5659GAT_2157_gat) );
AND2XL U_g2127 (.A(G1116GAT_96_ngat), .B(G5587GAT_2114_ngat), .Y(G5654GAT_2158_gat) );
AND2XL U_g2128 (.A(G921GAT_161_ngat), .B(G5569GAT_2131_ngat), .Y(G5638GAT_2159_gat) );
AND2XL U_g2129 (.A(G873GAT_177_ngat), .B(G5566GAT_2121_ngat), .Y(G5633GAT_2160_gat) );
AND2XL U_g2130 (.A(G5548GAT_2133_ngat), .B(G5374GAT_2056_ngat), .Y(G5618GAT_2161_gat) );
AND2XL U_g2131 (.A(G678GAT_242_ngat), .B(G5548GAT_2133_ngat), .Y(G5617GAT_2162_gat) );
AND2XL U_g2132 (.A(G5544GAT_2134_ngat), .B(G5370GAT_2057_ngat), .Y(G5613GAT_2163_gat) );
AND2XL U_g2133 (.A(G630GAT_258_ngat), .B(G5544GAT_2134_ngat), .Y(G5612GAT_2164_gat) );
AND2XL U_g2134 (.A(G5540GAT_2135_ngat), .B(G5366GAT_2058_ngat), .Y(G5608GAT_2165_gat) );
AND2XL U_g2135 (.A(G582GAT_274_ngat), .B(G5540GAT_2135_ngat), .Y(G5607GAT_2166_gat) );
AND2XL U_g2136 (.A(G5671GAT_2137_ngat), .B(G5670GAT_2136_ngat), .Y(G5727GAT_2167_gat) );
AND2XL U_g2137 (.A(G5666GAT_2138_ngat), .B(G5599GAT_2111_ngat), .Y(G5725GAT_2168_gat) );
AND2XL U_g2138 (.A(G5596GAT_2112_ngat), .B(G5666GAT_2138_ngat), .Y(G5726GAT_2169_gat) );
AND2XL U_g2139 (.A(G5660GAT_2140_ngat), .B(G5663GAT_2139_ngat), .Y(G5721GAT_2170_gat) );
AND2XL U_g2140 (.A(G5659GAT_2157_ngat), .B(G5658GAT_2141_ngat), .Y(G5718GAT_2171_gat) );
AND2XL U_g2141 (.A(G5654GAT_2158_ngat), .B(G5467GAT_2062_ngat), .Y(G5715GAT_2172_gat) );
AND2XL U_g2142 (.A(G5654GAT_2158_ngat), .B(G5587GAT_2114_ngat), .Y(G5713GAT_2173_gat) );
AND2XL U_g2143 (.A(G5650GAT_2144_ngat), .B(G5649GAT_2143_ngat), .Y(G5706GAT_2174_gat) );
AND2XL U_g2144 (.A(G5645GAT_2145_ngat), .B(G5578GAT_2118_ngat), .Y(G5704GAT_2175_gat) );
AND2XL U_g2145 (.A(G5575GAT_2119_ngat), .B(G5645GAT_2145_ngat), .Y(G5705GAT_2176_gat) );
AND2XL U_g2146 (.A(G5639GAT_2147_ngat), .B(G5642GAT_2146_ngat), .Y(G5700GAT_2177_gat) );
AND2XL U_g2147 (.A(G5638GAT_2159_ngat), .B(G5637GAT_2148_ngat), .Y(G5697GAT_2178_gat) );
AND2XL U_g2148 (.A(G5633GAT_2160_ngat), .B(G5446GAT_2069_ngat), .Y(G5694GAT_2179_gat) );
AND2XL U_g2149 (.A(G5633GAT_2160_ngat), .B(G5566GAT_2121_ngat), .Y(G5692GAT_2180_gat) );
AND2XL U_g2150 (.A(G5629GAT_2151_ngat), .B(G5628GAT_2150_ngat), .Y(G5685GAT_2181_gat) );
AND2XL U_g2151 (.A(G5624GAT_2152_ngat), .B(G5557GAT_2125_ngat), .Y(G5683GAT_2182_gat) );
AND2XL U_g2152 (.A(G5554GAT_2126_ngat), .B(G5624GAT_2152_ngat), .Y(G5684GAT_2183_gat) );
AND2XL U_g2153 (.A(G5618GAT_2161_ngat), .B(G5621GAT_2153_ngat), .Y(G5679GAT_2184_gat) );
AND2XL U_g2154 (.A(G5617GAT_2162_ngat), .B(G5616GAT_2154_ngat), .Y(G5676GAT_2185_gat) );
AND2XL U_g2155 (.A(G5612GAT_2164_ngat), .B(G5611GAT_2155_ngat), .Y(G5673GAT_2186_gat) );
AND2XL U_g2156 (.A(G5607GAT_2166_ngat), .B(G5606GAT_2156_ngat), .Y(G5672GAT_2187_gat) );
AND2XL U_g2157 (.A(G1116GAT_96_ngat), .B(G5654GAT_2158_ngat), .Y(G5714GAT_2188_gat) );
AND2XL U_g2158 (.A(G1068GAT_112_ngat), .B(G5651GAT_2142_ngat), .Y(G5709GAT_2189_gat) );
AND2XL U_g2159 (.A(G873GAT_177_ngat), .B(G5633GAT_2160_ngat), .Y(G5693GAT_2190_gat) );
AND2XL U_g2160 (.A(G825GAT_193_ngat), .B(G5630GAT_2149_ngat), .Y(G5688GAT_2191_gat) );
AND2XL U_g2161 (.A(G5726GAT_2169_ngat), .B(G5725GAT_2168_ngat), .Y(G5782GAT_2192_gat) );
AND2XL U_g2162 (.A(G5721GAT_2170_ngat), .B(G5663GAT_2139_ngat), .Y(G5780GAT_2193_gat) );
AND2XL U_g2163 (.A(G5660GAT_2140_ngat), .B(G5721GAT_2170_ngat), .Y(G5781GAT_2194_gat) );
AND2XL U_g2164 (.A(G5715GAT_2172_ngat), .B(G5718GAT_2171_ngat), .Y(G5776GAT_2195_gat) );
AND2XL U_g2165 (.A(G5714GAT_2188_ngat), .B(G5713GAT_2173_ngat), .Y(G5773GAT_2196_gat) );
AND2XL U_g2166 (.A(G5709GAT_2189_ngat), .B(G5522GAT_2090_ngat), .Y(G5770GAT_2197_gat) );
AND2XL U_g2167 (.A(G5709GAT_2189_ngat), .B(G5651GAT_2142_ngat), .Y(G5768GAT_2198_gat) );
AND2XL U_g2168 (.A(G5705GAT_2176_ngat), .B(G5704GAT_2175_ngat), .Y(G5761GAT_2199_gat) );
AND2XL U_g2169 (.A(G5700GAT_2177_ngat), .B(G5642GAT_2146_ngat), .Y(G5759GAT_2200_gat) );
AND2XL U_g2170 (.A(G5639GAT_2147_ngat), .B(G5700GAT_2177_ngat), .Y(G5760GAT_2201_gat) );
AND2XL U_g2171 (.A(G5694GAT_2179_ngat), .B(G5697GAT_2178_ngat), .Y(G5755GAT_2202_gat) );
AND2XL U_g2172 (.A(G5693GAT_2190_ngat), .B(G5692GAT_2180_ngat), .Y(G5752GAT_2203_gat) );
AND2XL U_g2173 (.A(G5688GAT_2191_ngat), .B(G5501GAT_2097_ngat), .Y(G5749GAT_2204_gat) );
AND2XL U_g2174 (.A(G5688GAT_2191_ngat), .B(G5630GAT_2149_ngat), .Y(G5747GAT_2205_gat) );
AND2XL U_g2175 (.A(G5684GAT_2183_ngat), .B(G5683GAT_2182_ngat), .Y(G5740GAT_2206_gat) );
AND2XL U_g2176 (.A(G5679GAT_2184_ngat), .B(G5621GAT_2153_ngat), .Y(G5738GAT_2207_gat) );
AND2XL U_g2177 (.A(G1068GAT_112_ngat), .B(G5709GAT_2189_ngat), .Y(G5769GAT_2208_gat) );
AND2XL U_g2178 (.A(G1020GAT_128_ngat), .B(G5706GAT_2174_ngat), .Y(G5764GAT_2209_gat) );
AND2XL U_g2179 (.A(G825GAT_193_ngat), .B(G5688GAT_2191_ngat), .Y(G5748GAT_2210_gat) );
AND2XL U_g2180 (.A(G777GAT_209_ngat), .B(G5685GAT_2181_ngat), .Y(G5743GAT_2211_gat) );
AND2XL U_g2181 (.A(G5618GAT_2161_ngat), .B(G5679GAT_2184_ngat), .Y(G5739GAT_2212_gat) );
AND2XL U_g2182 (.A(G5613GAT_2163_ngat), .B(G5676GAT_2185_ngat), .Y(G5734GAT_2213_gat) );
AND2XL U_g2183 (.A(G5608GAT_2165_ngat), .B(G5673GAT_2186_ngat), .Y(G5730GAT_2214_gat) );
AND2XL U_g2184 (.A(G5781GAT_2194_ngat), .B(G5780GAT_2193_ngat), .Y(G5831GAT_2215_gat) );
AND2XL U_g2185 (.A(G5776GAT_2195_ngat), .B(G5718GAT_2171_ngat), .Y(G5829GAT_2216_gat) );
AND2XL U_g2186 (.A(G5715GAT_2172_ngat), .B(G5776GAT_2195_ngat), .Y(G5830GAT_2217_gat) );
AND2XL U_g2187 (.A(G5770GAT_2197_ngat), .B(G5773GAT_2196_ngat), .Y(G5825GAT_2218_gat) );
AND2XL U_g2188 (.A(G5769GAT_2208_ngat), .B(G5768GAT_2198_ngat), .Y(G5822GAT_2219_gat) );
AND2XL U_g2189 (.A(G5764GAT_2209_ngat), .B(G5581GAT_2117_ngat), .Y(G5819GAT_2220_gat) );
AND2XL U_g2190 (.A(G5764GAT_2209_ngat), .B(G5706GAT_2174_ngat), .Y(G5817GAT_2221_gat) );
AND2XL U_g2191 (.A(G5760GAT_2201_ngat), .B(G5759GAT_2200_ngat), .Y(G5810GAT_2222_gat) );
AND2XL U_g2192 (.A(G5755GAT_2202_ngat), .B(G5697GAT_2178_ngat), .Y(G5808GAT_2223_gat) );
AND2XL U_g2193 (.A(G5694GAT_2179_ngat), .B(G5755GAT_2202_ngat), .Y(G5809GAT_2224_gat) );
AND2XL U_g2194 (.A(G5749GAT_2204_ngat), .B(G5752GAT_2203_ngat), .Y(G5804GAT_2225_gat) );
AND2XL U_g2195 (.A(G5748GAT_2210_ngat), .B(G5747GAT_2205_ngat), .Y(G5801GAT_2226_gat) );
AND2XL U_g2196 (.A(G5743GAT_2211_ngat), .B(G5560GAT_2124_ngat), .Y(G5798GAT_2227_gat) );
AND2XL U_g2197 (.A(G5743GAT_2211_ngat), .B(G5685GAT_2181_ngat), .Y(G5796GAT_2228_gat) );
AND2XL U_g2198 (.A(G5739GAT_2212_ngat), .B(G5738GAT_2207_ngat), .Y(G5789GAT_2229_gat) );
AND2XL U_g2199 (.A(G5734GAT_2213_ngat), .B(G5676GAT_2185_ngat), .Y(G5787GAT_2230_gat) );
AND2XL U_g2200 (.A(G5730GAT_2214_ngat), .B(G5673GAT_2186_ngat), .Y(G5785GAT_2231_gat) );
AND2XL U_g2201 (.A(G1020GAT_128_ngat), .B(G5764GAT_2209_ngat), .Y(G5818GAT_2232_gat) );
AND2XL U_g2202 (.A(G972GAT_144_ngat), .B(G5761GAT_2199_ngat), .Y(G5813GAT_2233_gat) );
AND2XL U_g2203 (.A(G777GAT_209_ngat), .B(G5743GAT_2211_ngat), .Y(G5797GAT_2234_gat) );
AND2XL U_g2204 (.A(G729GAT_225_ngat), .B(G5740GAT_2206_ngat), .Y(G5792GAT_2235_gat) );
AND2XL U_g2205 (.A(G5613GAT_2163_ngat), .B(G5734GAT_2213_ngat), .Y(G5788GAT_2236_gat) );
AND2XL U_g2206 (.A(G5608GAT_2165_ngat), .B(G5730GAT_2214_ngat), .Y(G5786GAT_2237_gat) );
AND2XL U_g2207 (.A(G5830GAT_2217_ngat), .B(G5829GAT_2216_ngat), .Y(G5879GAT_2238_gat) );
AND2XL U_g2208 (.A(G5825GAT_2218_ngat), .B(G5773GAT_2196_ngat), .Y(G5877GAT_2239_gat) );
AND2XL U_g2209 (.A(G5770GAT_2197_ngat), .B(G5825GAT_2218_ngat), .Y(G5878GAT_2240_gat) );
AND2XL U_g2210 (.A(G5819GAT_2220_ngat), .B(G5822GAT_2219_ngat), .Y(G5873GAT_2241_gat) );
AND2XL U_g2211 (.A(G5818GAT_2232_ngat), .B(G5817GAT_2221_ngat), .Y(G5870GAT_2242_gat) );
AND2XL U_g2212 (.A(G5813GAT_2233_ngat), .B(G5645GAT_2145_ngat), .Y(G5867GAT_2243_gat) );
AND2XL U_g2213 (.A(G5813GAT_2233_ngat), .B(G5761GAT_2199_ngat), .Y(G5865GAT_2244_gat) );
AND2XL U_g2214 (.A(G5809GAT_2224_ngat), .B(G5808GAT_2223_ngat), .Y(G5858GAT_2245_gat) );
AND2XL U_g2215 (.A(G5804GAT_2225_ngat), .B(G5752GAT_2203_ngat), .Y(G5856GAT_2246_gat) );
AND2XL U_g2216 (.A(G5749GAT_2204_ngat), .B(G5804GAT_2225_ngat), .Y(G5857GAT_2247_gat) );
AND2XL U_g2217 (.A(G5798GAT_2227_ngat), .B(G5801GAT_2226_ngat), .Y(G5852GAT_2248_gat) );
AND2XL U_g2218 (.A(G5797GAT_2234_ngat), .B(G5796GAT_2228_ngat), .Y(G5849GAT_2249_gat) );
AND2XL U_g2219 (.A(G5792GAT_2235_ngat), .B(G5624GAT_2152_ngat), .Y(G5846GAT_2250_gat) );
AND2XL U_g2220 (.A(G5792GAT_2235_ngat), .B(G5740GAT_2206_ngat), .Y(G5844GAT_2251_gat) );
AND2XL U_g2221 (.A(G5788GAT_2236_ngat), .B(G5787GAT_2230_ngat), .Y(G5837GAT_2252_gat) );
AND2XL U_g2222 (.A(G5786GAT_2237_ngat), .B(G5785GAT_2231_ngat), .Y(G5834GAT_2253_gat) );
AND2XL U_g2223 (.A(G972GAT_144_ngat), .B(G5813GAT_2233_ngat), .Y(G5866GAT_2254_gat) );
AND2XL U_g2224 (.A(G924GAT_160_ngat), .B(G5810GAT_2222_ngat), .Y(G5861GAT_2255_gat) );
AND2XL U_g2225 (.A(G729GAT_225_ngat), .B(G5792GAT_2235_ngat), .Y(G5845GAT_2256_gat) );
AND2XL U_g2226 (.A(G681GAT_241_ngat), .B(G5789GAT_2229_ngat), .Y(G5840GAT_2257_gat) );
AND2XL U_g2227 (.A(G5878GAT_2240_ngat), .B(G5877GAT_2239_ngat), .Y(G5925GAT_2258_gat) );
AND2XL U_g2228 (.A(G5873GAT_2241_ngat), .B(G5822GAT_2219_ngat), .Y(G5923GAT_2259_gat) );
AND2XL U_g2229 (.A(G5819GAT_2220_ngat), .B(G5873GAT_2241_ngat), .Y(G5924GAT_2260_gat) );
AND2XL U_g2230 (.A(G5867GAT_2243_ngat), .B(G5870GAT_2242_ngat), .Y(G5919GAT_2261_gat) );
AND2XL U_g2231 (.A(G5866GAT_2254_ngat), .B(G5865GAT_2244_ngat), .Y(G5916GAT_2262_gat) );
AND2XL U_g2232 (.A(G5861GAT_2255_ngat), .B(G5700GAT_2177_ngat), .Y(G5913GAT_2263_gat) );
AND2XL U_g2233 (.A(G5861GAT_2255_ngat), .B(G5810GAT_2222_ngat), .Y(G5911GAT_2264_gat) );
AND2XL U_g2234 (.A(G5857GAT_2247_ngat), .B(G5856GAT_2246_ngat), .Y(G5904GAT_2265_gat) );
AND2XL U_g2235 (.A(G5852GAT_2248_ngat), .B(G5801GAT_2226_ngat), .Y(G5902GAT_2266_gat) );
AND2XL U_g2236 (.A(G5798GAT_2227_ngat), .B(G5852GAT_2248_ngat), .Y(G5903GAT_2267_gat) );
AND2XL U_g2237 (.A(G5846GAT_2250_ngat), .B(G5849GAT_2249_ngat), .Y(G5898GAT_2268_gat) );
AND2XL U_g2238 (.A(G5845GAT_2256_ngat), .B(G5844GAT_2251_ngat), .Y(G5895GAT_2269_gat) );
AND2XL U_g2239 (.A(G5840GAT_2257_ngat), .B(G5679GAT_2184_ngat), .Y(G5892GAT_2270_gat) );
AND2XL U_g2240 (.A(G5840GAT_2257_ngat), .B(G5789GAT_2229_ngat), .Y(G5890GAT_2271_gat) );
AND2XL U_g2241 (.A(G924GAT_160_ngat), .B(G5861GAT_2255_ngat), .Y(G5912GAT_2272_gat) );
AND2XL U_g2242 (.A(G876GAT_176_ngat), .B(G5858GAT_2245_ngat), .Y(G5907GAT_2273_gat) );
AND2XL U_g2243 (.A(G681GAT_241_ngat), .B(G5840GAT_2257_ngat), .Y(G5891GAT_2274_gat) );
AND2XL U_g2244 (.A(G633GAT_257_ngat), .B(G5837GAT_2252_ngat), .Y(G5886GAT_2275_gat) );
AND2XL U_g2245 (.A(G585GAT_273_ngat), .B(G5834GAT_2253_ngat), .Y(G5882GAT_2276_gat) );
AND2XL U_g2246 (.A(G5924GAT_2260_ngat), .B(G5923GAT_2259_ngat), .Y(G5968GAT_2277_gat) );
AND2XL U_g2247 (.A(G5919GAT_2261_ngat), .B(G5870GAT_2242_ngat), .Y(G5966GAT_2278_gat) );
AND2XL U_g2248 (.A(G5867GAT_2243_ngat), .B(G5919GAT_2261_ngat), .Y(G5967GAT_2279_gat) );
AND2XL U_g2249 (.A(G5913GAT_2263_ngat), .B(G5916GAT_2262_ngat), .Y(G5962GAT_2280_gat) );
AND2XL U_g2250 (.A(G5912GAT_2272_ngat), .B(G5911GAT_2264_ngat), .Y(G5959GAT_2281_gat) );
AND2XL U_g2251 (.A(G5907GAT_2273_ngat), .B(G5755GAT_2202_ngat), .Y(G5956GAT_2282_gat) );
AND2XL U_g2252 (.A(G5907GAT_2273_ngat), .B(G5858GAT_2245_ngat), .Y(G5954GAT_2283_gat) );
AND2XL U_g2253 (.A(G5903GAT_2267_ngat), .B(G5902GAT_2266_ngat), .Y(G5947GAT_2284_gat) );
AND2XL U_g2254 (.A(G5898GAT_2268_ngat), .B(G5849GAT_2249_ngat), .Y(G5945GAT_2285_gat) );
AND2XL U_g2255 (.A(G5846GAT_2250_ngat), .B(G5898GAT_2268_ngat), .Y(G5946GAT_2286_gat) );
AND2XL U_g2256 (.A(G5892GAT_2270_ngat), .B(G5895GAT_2269_ngat), .Y(G5941GAT_2287_gat) );
AND2XL U_g2257 (.A(G5891GAT_2274_ngat), .B(G5890GAT_2271_ngat), .Y(G5938GAT_2288_gat) );
AND2XL U_g2258 (.A(G5886GAT_2275_ngat), .B(G5837GAT_2252_ngat), .Y(G5933GAT_2289_gat) );
AND2XL U_g2259 (.A(G5882GAT_2276_ngat), .B(G5834GAT_2253_ngat), .Y(G5928GAT_2290_gat) );
AND2XL U_g2260 (.A(G876GAT_176_ngat), .B(G5907GAT_2273_ngat), .Y(G5955GAT_2291_gat) );
AND2XL U_g2261 (.A(G828GAT_192_ngat), .B(G5904GAT_2265_ngat), .Y(G5950GAT_2292_gat) );
AND2XL U_g2262 (.A(G5886GAT_2275_ngat), .B(G5734GAT_2213_ngat), .Y(G5935GAT_2293_gat) );
AND2XL U_g2263 (.A(G633GAT_257_ngat), .B(G5886GAT_2275_ngat), .Y(G5934GAT_2294_gat) );
AND2XL U_g2264 (.A(G5882GAT_2276_ngat), .B(G5730GAT_2214_ngat), .Y(G5930GAT_2295_gat) );
AND2XL U_g2265 (.A(G585GAT_273_ngat), .B(G5882GAT_2276_ngat), .Y(G5929GAT_2296_gat) );
AND2XL U_g2266 (.A(G5967GAT_2279_ngat), .B(G5966GAT_2278_ngat), .Y(G6002GAT_2297_gat) );
AND2XL U_g2267 (.A(G5962GAT_2280_ngat), .B(G5916GAT_2262_ngat), .Y(G6000GAT_2298_gat) );
AND2XL U_g2268 (.A(G5913GAT_2263_ngat), .B(G5962GAT_2280_ngat), .Y(G6001GAT_2299_gat) );
AND2XL U_g2269 (.A(G5956GAT_2282_ngat), .B(G5959GAT_2281_ngat), .Y(G5996GAT_2300_gat) );
AND2XL U_g2270 (.A(G5955GAT_2291_ngat), .B(G5954GAT_2283_ngat), .Y(G5993GAT_2301_gat) );
AND2XL U_g2271 (.A(G5950GAT_2292_ngat), .B(G5804GAT_2225_ngat), .Y(G5990GAT_2302_gat) );
AND2XL U_g2272 (.A(G5950GAT_2292_ngat), .B(G5904GAT_2265_ngat), .Y(G5988GAT_2303_gat) );
AND2XL U_g2273 (.A(G5946GAT_2286_ngat), .B(G5945GAT_2285_ngat), .Y(G5981GAT_2304_gat) );
AND2XL U_g2274 (.A(G5941GAT_2287_ngat), .B(G5895GAT_2269_ngat), .Y(G5979GAT_2305_gat) );
AND2XL U_g2275 (.A(G5892GAT_2270_ngat), .B(G5941GAT_2287_ngat), .Y(G5980GAT_2306_gat) );
AND2XL U_g2276 (.A(G5935GAT_2293_ngat), .B(G5938GAT_2288_ngat), .Y(G5975GAT_2307_gat) );
AND2XL U_g2277 (.A(G5934GAT_2294_ngat), .B(G5933GAT_2289_ngat), .Y(G5972GAT_2308_gat) );
AND2XL U_g2278 (.A(G5929GAT_2296_ngat), .B(G5928GAT_2290_ngat), .Y(G5971GAT_2309_gat) );
AND2XL U_g2279 (.A(G828GAT_192_ngat), .B(G5950GAT_2292_ngat), .Y(G5989GAT_2310_gat) );
AND2XL U_g2280 (.A(G780GAT_208_ngat), .B(G5947GAT_2284_ngat), .Y(G5984GAT_2311_gat) );
AND2XL U_g2281 (.A(G6001GAT_2299_ngat), .B(G6000GAT_2298_ngat), .Y(G6032GAT_2312_gat) );
AND2XL U_g2282 (.A(G5996GAT_2300_ngat), .B(G5959GAT_2281_ngat), .Y(G6030GAT_2313_gat) );
AND2XL U_g2283 (.A(G5956GAT_2282_ngat), .B(G5996GAT_2300_ngat), .Y(G6031GAT_2314_gat) );
AND2XL U_g2284 (.A(G5990GAT_2302_ngat), .B(G5993GAT_2301_ngat), .Y(G6026GAT_2315_gat) );
AND2XL U_g2285 (.A(G5989GAT_2310_ngat), .B(G5988GAT_2303_ngat), .Y(G6023GAT_2316_gat) );
AND2XL U_g2286 (.A(G5984GAT_2311_ngat), .B(G5852GAT_2248_ngat), .Y(G6020GAT_2317_gat) );
AND2XL U_g2287 (.A(G5984GAT_2311_ngat), .B(G5947GAT_2284_ngat), .Y(G6018GAT_2318_gat) );
AND2XL U_g2288 (.A(G5980GAT_2306_ngat), .B(G5979GAT_2305_ngat), .Y(G6011GAT_2319_gat) );
AND2XL U_g2289 (.A(G5975GAT_2307_ngat), .B(G5938GAT_2288_ngat), .Y(G6009GAT_2320_gat) );
AND2XL U_g2290 (.A(G780GAT_208_ngat), .B(G5984GAT_2311_ngat), .Y(G6019GAT_2321_gat) );
AND2XL U_g2291 (.A(G732GAT_224_ngat), .B(G5981GAT_2304_ngat), .Y(G6014GAT_2322_gat) );
AND2XL U_g2292 (.A(G5935GAT_2293_ngat), .B(G5975GAT_2307_ngat), .Y(G6010GAT_2323_gat) );
AND2XL U_g2293 (.A(G5930GAT_2295_ngat), .B(G5972GAT_2308_ngat), .Y(G6005GAT_2324_gat) );
AND2XL U_g2294 (.A(G6031GAT_2314_ngat), .B(G6030GAT_2313_ngat), .Y(G6058GAT_2325_gat) );
AND2XL U_g2295 (.A(G6026GAT_2315_ngat), .B(G5993GAT_2301_ngat), .Y(G6056GAT_2326_gat) );
AND2XL U_g2296 (.A(G5990GAT_2302_ngat), .B(G6026GAT_2315_ngat), .Y(G6057GAT_2327_gat) );
AND2XL U_g2297 (.A(G6020GAT_2317_ngat), .B(G6023GAT_2316_ngat), .Y(G6052GAT_2328_gat) );
AND2XL U_g2298 (.A(G6019GAT_2321_ngat), .B(G6018GAT_2318_ngat), .Y(G6049GAT_2329_gat) );
AND2XL U_g2299 (.A(G6014GAT_2322_ngat), .B(G5898GAT_2268_ngat), .Y(G6046GAT_2330_gat) );
AND2XL U_g2300 (.A(G6014GAT_2322_ngat), .B(G5981GAT_2304_ngat), .Y(G6044GAT_2331_gat) );
AND2XL U_g2301 (.A(G6010GAT_2323_ngat), .B(G6009GAT_2320_ngat), .Y(G6037GAT_2332_gat) );
AND2XL U_g2302 (.A(G6005GAT_2324_ngat), .B(G5972GAT_2308_ngat), .Y(G6035GAT_2333_gat) );
AND2XL U_g2303 (.A(G732GAT_224_ngat), .B(G6014GAT_2322_ngat), .Y(G6045GAT_2334_gat) );
AND2XL U_g2304 (.A(G684GAT_240_ngat), .B(G6011GAT_2319_ngat), .Y(G6040GAT_2335_gat) );
AND2XL U_g2305 (.A(G5930GAT_2295_ngat), .B(G6005GAT_2324_ngat), .Y(G6036GAT_2336_gat) );
AND2XL U_g2306 (.A(G6057GAT_2327_ngat), .B(G6056GAT_2326_ngat), .Y(G6082GAT_2337_gat) );
AND2XL U_g2307 (.A(G6052GAT_2328_ngat), .B(G6023GAT_2316_ngat), .Y(G6080GAT_2338_gat) );
AND2XL U_g2308 (.A(G6020GAT_2317_ngat), .B(G6052GAT_2328_ngat), .Y(G6081GAT_2339_gat) );
AND2XL U_g2309 (.A(G6046GAT_2330_ngat), .B(G6049GAT_2329_ngat), .Y(G6076GAT_2340_gat) );
AND2XL U_g2310 (.A(G6045GAT_2334_ngat), .B(G6044GAT_2331_ngat), .Y(G6073GAT_2341_gat) );
AND2XL U_g2311 (.A(G6040GAT_2335_ngat), .B(G5941GAT_2287_ngat), .Y(G6070GAT_2342_gat) );
AND2XL U_g2312 (.A(G6040GAT_2335_ngat), .B(G6011GAT_2319_ngat), .Y(G6068GAT_2343_gat) );
AND2XL U_g2313 (.A(G6036GAT_2336_ngat), .B(G6035GAT_2333_ngat), .Y(G6061GAT_2344_gat) );
AND2XL U_g2314 (.A(G684GAT_240_ngat), .B(G6040GAT_2335_ngat), .Y(G6069GAT_2345_gat) );
AND2XL U_g2315 (.A(G636GAT_256_ngat), .B(G6037GAT_2332_ngat), .Y(G6064GAT_2346_gat) );
AND2XL U_g2316 (.A(G6081GAT_2339_ngat), .B(G6080GAT_2338_ngat), .Y(G6103GAT_2347_gat) );
AND2XL U_g2317 (.A(G6076GAT_2340_ngat), .B(G6049GAT_2329_ngat), .Y(G6101GAT_2348_gat) );
AND2XL U_g2318 (.A(G6046GAT_2330_ngat), .B(G6076GAT_2340_ngat), .Y(G6102GAT_2349_gat) );
AND2XL U_g2319 (.A(G6070GAT_2342_ngat), .B(G6073GAT_2341_ngat), .Y(G6097GAT_2350_gat) );
AND2XL U_g2320 (.A(G6069GAT_2345_ngat), .B(G6068GAT_2343_ngat), .Y(G6094GAT_2351_gat) );
AND2XL U_g2321 (.A(G6064GAT_2346_ngat), .B(G5975GAT_2307_ngat), .Y(G6091GAT_2352_gat) );
AND2XL U_g2322 (.A(G6064GAT_2346_ngat), .B(G6037GAT_2332_ngat), .Y(G6089GAT_2353_gat) );
AND2XL U_g2323 (.A(G636GAT_256_ngat), .B(G6064GAT_2346_ngat), .Y(G6090GAT_2354_gat) );
AND2XL U_g2324 (.A(G588GAT_272_ngat), .B(G6061GAT_2344_ngat), .Y(G6085GAT_2355_gat) );
AND2XL U_g2325 (.A(G6102GAT_2349_ngat), .B(G6101GAT_2348_ngat), .Y(G6120GAT_2356_gat) );
AND2XL U_g2326 (.A(G6097GAT_2350_ngat), .B(G6073GAT_2341_ngat), .Y(G6118GAT_2357_gat) );
AND2XL U_g2327 (.A(G6070GAT_2342_ngat), .B(G6097GAT_2350_ngat), .Y(G6119GAT_2358_gat) );
AND2XL U_g2328 (.A(G6091GAT_2352_ngat), .B(G6094GAT_2351_ngat), .Y(G6114GAT_2359_gat) );
AND2XL U_g2329 (.A(G6090GAT_2354_ngat), .B(G6089GAT_2353_ngat), .Y(G6111GAT_2360_gat) );
AND2XL U_g2330 (.A(G6085GAT_2355_ngat), .B(G6061GAT_2344_ngat), .Y(G6106GAT_2361_gat) );
AND2XL U_g2331 (.A(G6085GAT_2355_ngat), .B(G6005GAT_2324_ngat), .Y(G6108GAT_2362_gat) );
AND2XL U_g2332 (.A(G588GAT_272_ngat), .B(G6085GAT_2355_ngat), .Y(G6107GAT_2363_gat) );
AND2XL U_g2333 (.A(G6119GAT_2358_ngat), .B(G6118GAT_2357_ngat), .Y(G6130GAT_2364_gat) );
AND2XL U_g2334 (.A(G6114GAT_2359_ngat), .B(G6094GAT_2351_ngat), .Y(G6128GAT_2365_gat) );
AND2XL U_g2335 (.A(G6091GAT_2352_ngat), .B(G6114GAT_2359_ngat), .Y(G6129GAT_2366_gat) );
AND2XL U_g2336 (.A(G6108GAT_2362_ngat), .B(G6111GAT_2360_ngat), .Y(G6124GAT_2367_gat) );
AND2XL U_g2337 (.A(G6107GAT_2363_ngat), .B(G6106GAT_2361_ngat), .Y(G6123GAT_2368_gat) );
AND2XL U_g2338 (.A(G6129GAT_2366_ngat), .B(G6128GAT_2365_ngat), .Y(G6135GAT_2369_gat) );
AND2XL U_g2339 (.A(G6124GAT_2367_ngat), .B(G6111GAT_2360_ngat), .Y(G6133GAT_2370_gat) );
AND2XL U_g2340 (.A(G6108GAT_2362_ngat), .B(G6124GAT_2367_ngat), .Y(G6134GAT_2371_gat) );
AND2XL U_g2341 (.A(G6134GAT_2371_ngat), .B(G6133GAT_2370_ngat), .Y(G6138GAT_2372_gat) );
BUFX20 U_g2342 (.A(G6138GAT_2372_gat), .Y(G6141GAT_2373_gat) );
AND2XL U_g2343 (.A(G6141GAT_2373_ngat), .B(G6124GAT_2367_ngat), .Y(G6147GAT_2374_gat) );
AND2XL U_g2344 (.A(G6141GAT_2373_ngat), .B(G6138GAT_2372_ngat), .Y(G6145GAT_2375_gat) );
BUFX20 U_g2345 (.A(G6141GAT_2373_gat), .Y(G6146GAT_2376_gat) );
AND2XL U_g2346 (.A(G6147GAT_2374_ngat), .B(G6135GAT_2369_ngat), .Y(G6151GAT_2377_gat) );
AND2XL U_g2347 (.A(G6146GAT_2376_ngat), .B(G6145GAT_2375_ngat), .Y(G6150GAT_2378_gat) );
AND2XL U_g2348 (.A(G6151GAT_2377_ngat), .B(G6114GAT_2359_ngat), .Y(G6157GAT_2379_gat) );
AND2XL U_g2349 (.A(G6151GAT_2377_ngat), .B(G6135GAT_2369_ngat), .Y(G6155GAT_2380_gat) );
AND2XL U_g2350 (.A(G6147GAT_2374_ngat), .B(G6151GAT_2377_ngat), .Y(G6156GAT_2381_gat) );
AND2XL U_g2351 (.A(G6157GAT_2379_ngat), .B(G6130GAT_2364_ngat), .Y(G6161GAT_2382_gat) );
AND2XL U_g2352 (.A(G6156GAT_2381_ngat), .B(G6155GAT_2380_ngat), .Y(G6160GAT_2383_gat) );
AND2XL U_g2353 (.A(G6161GAT_2382_ngat), .B(G6097GAT_2350_ngat), .Y(G6167GAT_2384_gat) );
AND2XL U_g2354 (.A(G6161GAT_2382_ngat), .B(G6130GAT_2364_ngat), .Y(G6165GAT_2385_gat) );
AND2XL U_g2355 (.A(G6157GAT_2379_ngat), .B(G6161GAT_2382_ngat), .Y(G6166GAT_2386_gat) );
AND2XL U_g2356 (.A(G6167GAT_2384_ngat), .B(G6120GAT_2356_ngat), .Y(G6171GAT_2387_gat) );
AND2XL U_g2357 (.A(G6166GAT_2386_ngat), .B(G6165GAT_2385_ngat), .Y(G6170GAT_2388_gat) );
AND2XL U_g2358 (.A(G6171GAT_2387_ngat), .B(G6076GAT_2340_ngat), .Y(G6177GAT_2389_gat) );
AND2XL U_g2359 (.A(G6171GAT_2387_ngat), .B(G6120GAT_2356_ngat), .Y(G6175GAT_2390_gat) );
AND2XL U_g2360 (.A(G6167GAT_2384_ngat), .B(G6171GAT_2387_ngat), .Y(G6176GAT_2391_gat) );
AND2XL U_g2361 (.A(G6177GAT_2389_ngat), .B(G6103GAT_2347_ngat), .Y(G6181GAT_2392_gat) );
AND2XL U_g2362 (.A(G6176GAT_2391_ngat), .B(G6175GAT_2390_ngat), .Y(G6180GAT_2393_gat) );
AND2XL U_g2363 (.A(G6181GAT_2392_ngat), .B(G6052GAT_2328_ngat), .Y(G6187GAT_2394_gat) );
AND2XL U_g2364 (.A(G6181GAT_2392_ngat), .B(G6103GAT_2347_ngat), .Y(G6185GAT_2395_gat) );
AND2XL U_g2365 (.A(G6177GAT_2389_ngat), .B(G6181GAT_2392_ngat), .Y(G6186GAT_2396_gat) );
AND2XL U_g2366 (.A(G6187GAT_2394_ngat), .B(G6082GAT_2337_ngat), .Y(G6191GAT_2397_gat) );
AND2XL U_g2367 (.A(G6186GAT_2396_ngat), .B(G6185GAT_2395_ngat), .Y(G6190GAT_2398_gat) );
AND2XL U_g2368 (.A(G6191GAT_2397_ngat), .B(G6026GAT_2315_ngat), .Y(G6197GAT_2399_gat) );
AND2XL U_g2369 (.A(G6191GAT_2397_ngat), .B(G6082GAT_2337_ngat), .Y(G6195GAT_2400_gat) );
AND2XL U_g2370 (.A(G6187GAT_2394_ngat), .B(G6191GAT_2397_ngat), .Y(G6196GAT_2401_gat) );
AND2XL U_g2371 (.A(G6197GAT_2399_ngat), .B(G6058GAT_2325_ngat), .Y(G6201GAT_2402_gat) );
AND2XL U_g2372 (.A(G6196GAT_2401_ngat), .B(G6195GAT_2400_ngat), .Y(G6200GAT_2403_gat) );
AND2XL U_g2373 (.A(G6201GAT_2402_ngat), .B(G5996GAT_2300_ngat), .Y(G6207GAT_2404_gat) );
AND2XL U_g2374 (.A(G6201GAT_2402_ngat), .B(G6058GAT_2325_ngat), .Y(G6205GAT_2405_gat) );
AND2XL U_g2375 (.A(G6197GAT_2399_ngat), .B(G6201GAT_2402_ngat), .Y(G6206GAT_2406_gat) );
AND2XL U_g2376 (.A(G6207GAT_2404_ngat), .B(G6032GAT_2312_ngat), .Y(G6211GAT_2407_gat) );
AND2XL U_g2377 (.A(G6206GAT_2406_ngat), .B(G6205GAT_2405_ngat), .Y(G6210GAT_2408_gat) );
AND2XL U_g2378 (.A(G6211GAT_2407_ngat), .B(G5962GAT_2280_ngat), .Y(G6217GAT_2409_gat) );
AND2XL U_g2379 (.A(G6211GAT_2407_ngat), .B(G6032GAT_2312_ngat), .Y(G6215GAT_2410_gat) );
AND2XL U_g2380 (.A(G6207GAT_2404_ngat), .B(G6211GAT_2407_ngat), .Y(G6216GAT_2411_gat) );
AND2XL U_g2381 (.A(G6217GAT_2409_ngat), .B(G6002GAT_2297_ngat), .Y(G6221GAT_2412_gat) );
AND2XL U_g2382 (.A(G6216GAT_2411_ngat), .B(G6215GAT_2410_ngat), .Y(G6220GAT_2413_gat) );
AND2XL U_g2383 (.A(G6221GAT_2412_ngat), .B(G5919GAT_2261_ngat), .Y(G6227GAT_2414_gat) );
AND2XL U_g2384 (.A(G6221GAT_2412_ngat), .B(G6002GAT_2297_ngat), .Y(G6225GAT_2415_gat) );
AND2XL U_g2385 (.A(G6217GAT_2409_ngat), .B(G6221GAT_2412_ngat), .Y(G6226GAT_2416_gat) );
AND2XL U_g2386 (.A(G6227GAT_2414_ngat), .B(G5968GAT_2277_ngat), .Y(G6231GAT_2417_gat) );
AND2XL U_g2387 (.A(G6226GAT_2416_ngat), .B(G6225GAT_2415_ngat), .Y(G6230GAT_2418_gat) );
AND2XL U_g2388 (.A(G6231GAT_2417_ngat), .B(G5873GAT_2241_ngat), .Y(G6237GAT_2419_gat) );
AND2XL U_g2389 (.A(G6231GAT_2417_ngat), .B(G5968GAT_2277_ngat), .Y(G6235GAT_2420_gat) );
AND2XL U_g2390 (.A(G6227GAT_2414_ngat), .B(G6231GAT_2417_ngat), .Y(G6236GAT_2421_gat) );
AND2XL U_g2391 (.A(G6237GAT_2419_ngat), .B(G5925GAT_2258_ngat), .Y(G6241GAT_2422_gat) );
AND2XL U_g2392 (.A(G6236GAT_2421_ngat), .B(G6235GAT_2420_ngat), .Y(G6240GAT_2423_gat) );
AND2XL U_g2393 (.A(G6241GAT_2422_ngat), .B(G5825GAT_2218_ngat), .Y(G6247GAT_2424_gat) );
AND2XL U_g2394 (.A(G6241GAT_2422_ngat), .B(G5925GAT_2258_ngat), .Y(G6245GAT_2425_gat) );
AND2XL U_g2395 (.A(G6237GAT_2419_ngat), .B(G6241GAT_2422_ngat), .Y(G6246GAT_2426_gat) );
AND2XL U_g2396 (.A(G6247GAT_2424_ngat), .B(G5879GAT_2238_ngat), .Y(G6251GAT_2427_gat) );
AND2XL U_g2397 (.A(G6246GAT_2426_ngat), .B(G6245GAT_2425_ngat), .Y(G6250GAT_2428_gat) );
AND2XL U_g2398 (.A(G6251GAT_2427_ngat), .B(G5776GAT_2195_ngat), .Y(G6257GAT_2429_gat) );
AND2XL U_g2399 (.A(G6251GAT_2427_ngat), .B(G5879GAT_2238_ngat), .Y(G6255GAT_2430_gat) );
AND2XL U_g2400 (.A(G6247GAT_2424_ngat), .B(G6251GAT_2427_ngat), .Y(G6256GAT_2431_gat) );
AND2XL U_g2401 (.A(G6257GAT_2429_ngat), .B(G5831GAT_2215_ngat), .Y(G6261GAT_2432_gat) );
AND2XL U_g2402 (.A(G6256GAT_2431_ngat), .B(G6255GAT_2430_ngat), .Y(G6260GAT_2433_gat) );
AND2XL U_g2403 (.A(G6261GAT_2432_ngat), .B(G5721GAT_2170_ngat), .Y(G6267GAT_2434_gat) );
AND2XL U_g2404 (.A(G6261GAT_2432_ngat), .B(G5831GAT_2215_ngat), .Y(G6265GAT_2435_gat) );
AND2XL U_g2405 (.A(G6257GAT_2429_ngat), .B(G6261GAT_2432_ngat), .Y(G6266GAT_2436_gat) );
AND2XL U_g2406 (.A(G6267GAT_2434_ngat), .B(G5782GAT_2192_ngat), .Y(G6271GAT_2437_gat) );
AND2XL U_g2407 (.A(G6266GAT_2436_ngat), .B(G6265GAT_2435_ngat), .Y(G6270GAT_2438_gat) );
AND2XL U_g2408 (.A(G6271GAT_2437_ngat), .B(G5666GAT_2138_ngat), .Y(G6277GAT_2439_gat) );
AND2XL U_g2409 (.A(G6271GAT_2437_ngat), .B(G5782GAT_2192_ngat), .Y(G6275GAT_2440_gat) );
AND2XL U_g2410 (.A(G6267GAT_2434_ngat), .B(G6271GAT_2437_ngat), .Y(G6276GAT_2441_gat) );
AND2XL U_g2411 (.A(G6277GAT_2439_ngat), .B(G5727GAT_2167_ngat), .Y(G6281GAT_2442_gat) );
AND2XL U_g2412 (.A(G6276GAT_2441_ngat), .B(G6275GAT_2440_ngat), .Y(G6280GAT_2443_gat) );
AND2XL U_g2413 (.A(G6281GAT_2442_ngat), .B(G5602GAT_2110_ngat), .Y(G6287GAT_2444_gat) );
AND2XL U_g2414 (.A(G6281GAT_2442_ngat), .B(G5727GAT_2167_ngat), .Y(G6285GAT_2445_gat) );
AND2XL U_g2415 (.A(G6277GAT_2439_ngat), .B(G6281GAT_2442_ngat), .Y(G6286GAT_2446_gat) );
AND2XL U_g2416 (.A(G6286GAT_2446_ngat), .B(G6285GAT_2445_ngat), .Y(G6288GAT_2447_gat) );
INVXL U_g2417 (.A(G1263GAT_47_gat), .Y(G1263GAT_47_ngat) );
INVXL U_g2418 (.A(G1367GAT_288_gat), .Y(G1367GAT_288_ngat) );
INVXL U_g2419 (.A(G1215GAT_63_gat), .Y(G1215GAT_63_ngat) );
INVXL U_g2420 (.A(G1363GAT_289_gat), .Y(G1363GAT_289_ngat) );
INVXL U_g2421 (.A(G1167GAT_79_gat), .Y(G1167GAT_79_ngat) );
INVXL U_g2422 (.A(G1359GAT_290_gat), .Y(G1359GAT_290_ngat) );
INVXL U_g2423 (.A(G1119GAT_95_gat), .Y(G1119GAT_95_ngat) );
INVXL U_g2424 (.A(G1355GAT_291_gat), .Y(G1355GAT_291_ngat) );
INVXL U_g2425 (.A(G1071GAT_111_gat), .Y(G1071GAT_111_ngat) );
INVXL U_g2426 (.A(G1351GAT_292_gat), .Y(G1351GAT_292_ngat) );
INVXL U_g2427 (.A(G1023GAT_127_gat), .Y(G1023GAT_127_ngat) );
INVXL U_g2428 (.A(G1347GAT_293_gat), .Y(G1347GAT_293_ngat) );
INVXL U_g2429 (.A(G975GAT_143_gat), .Y(G975GAT_143_ngat) );
INVXL U_g2430 (.A(G1343GAT_294_gat), .Y(G1343GAT_294_ngat) );
INVXL U_g2431 (.A(G927GAT_159_gat), .Y(G927GAT_159_ngat) );
INVXL U_g2432 (.A(G1339GAT_295_gat), .Y(G1339GAT_295_ngat) );
INVXL U_g2433 (.A(G879GAT_175_gat), .Y(G879GAT_175_ngat) );
INVXL U_g2434 (.A(G1335GAT_296_gat), .Y(G1335GAT_296_ngat) );
INVXL U_g2435 (.A(G831GAT_191_gat), .Y(G831GAT_191_ngat) );
INVXL U_g2436 (.A(G1331GAT_297_gat), .Y(G1331GAT_297_ngat) );
INVXL U_g2437 (.A(G783GAT_207_gat), .Y(G783GAT_207_ngat) );
INVXL U_g2438 (.A(G1327GAT_298_gat), .Y(G1327GAT_298_ngat) );
INVXL U_g2439 (.A(G735GAT_223_gat), .Y(G735GAT_223_ngat) );
INVXL U_g2440 (.A(G1323GAT_299_gat), .Y(G1323GAT_299_ngat) );
INVXL U_g2441 (.A(G687GAT_239_gat), .Y(G687GAT_239_ngat) );
INVXL U_g2442 (.A(G1319GAT_300_gat), .Y(G1319GAT_300_ngat) );
INVXL U_g2443 (.A(G639GAT_255_gat), .Y(G639GAT_255_ngat) );
INVXL U_g2444 (.A(G1315GAT_301_gat), .Y(G1315GAT_301_ngat) );
INVXL U_g2445 (.A(G591GAT_271_gat), .Y(G591GAT_271_ngat) );
INVXL U_g2446 (.A(G1311GAT_302_gat), .Y(G1311GAT_302_ngat) );
INVXL U_g2447 (.A(G1399GAT_304_gat), .Y(G1399GAT_304_ngat) );
INVXL U_g2448 (.A(G1400GAT_303_gat), .Y(G1400GAT_303_ngat) );
INVXL U_g2449 (.A(G1397GAT_306_gat), .Y(G1397GAT_306_ngat) );
INVXL U_g2450 (.A(G1398GAT_305_gat), .Y(G1398GAT_305_ngat) );
INVXL U_g2451 (.A(G1395GAT_308_gat), .Y(G1395GAT_308_ngat) );
INVXL U_g2452 (.A(G1396GAT_307_gat), .Y(G1396GAT_307_ngat) );
INVXL U_g2453 (.A(G1393GAT_310_gat), .Y(G1393GAT_310_ngat) );
INVXL U_g2454 (.A(G1394GAT_309_gat), .Y(G1394GAT_309_ngat) );
INVXL U_g2455 (.A(G1391GAT_312_gat), .Y(G1391GAT_312_ngat) );
INVXL U_g2456 (.A(G1392GAT_311_gat), .Y(G1392GAT_311_ngat) );
INVXL U_g2457 (.A(G1389GAT_314_gat), .Y(G1389GAT_314_ngat) );
INVXL U_g2458 (.A(G1390GAT_313_gat), .Y(G1390GAT_313_ngat) );
INVXL U_g2459 (.A(G1387GAT_316_gat), .Y(G1387GAT_316_ngat) );
INVXL U_g2460 (.A(G1388GAT_315_gat), .Y(G1388GAT_315_ngat) );
INVXL U_g2461 (.A(G1385GAT_318_gat), .Y(G1385GAT_318_ngat) );
INVXL U_g2462 (.A(G1386GAT_317_gat), .Y(G1386GAT_317_ngat) );
INVXL U_g2463 (.A(G1383GAT_320_gat), .Y(G1383GAT_320_ngat) );
INVXL U_g2464 (.A(G1384GAT_319_gat), .Y(G1384GAT_319_ngat) );
INVXL U_g2465 (.A(G1381GAT_322_gat), .Y(G1381GAT_322_ngat) );
INVXL U_g2466 (.A(G1382GAT_321_gat), .Y(G1382GAT_321_ngat) );
INVXL U_g2467 (.A(G1379GAT_324_gat), .Y(G1379GAT_324_ngat) );
INVXL U_g2468 (.A(G1380GAT_323_gat), .Y(G1380GAT_323_ngat) );
INVXL U_g2469 (.A(G1377GAT_326_gat), .Y(G1377GAT_326_ngat) );
INVXL U_g2470 (.A(G1378GAT_325_gat), .Y(G1378GAT_325_ngat) );
INVXL U_g2471 (.A(G1375GAT_328_gat), .Y(G1375GAT_328_ngat) );
INVXL U_g2472 (.A(G1376GAT_327_gat), .Y(G1376GAT_327_ngat) );
INVXL U_g2473 (.A(G1373GAT_330_gat), .Y(G1373GAT_330_ngat) );
INVXL U_g2474 (.A(G1374GAT_329_gat), .Y(G1374GAT_329_ngat) );
INVXL U_g2475 (.A(G1371GAT_332_gat), .Y(G1371GAT_332_ngat) );
INVXL U_g2476 (.A(G1372GAT_331_gat), .Y(G1372GAT_331_ngat) );
INVXL U_g2477 (.A(G1443GAT_333_gat), .Y(G1443GAT_333_ngat) );
INVXL U_g2478 (.A(G1218GAT_62_gat), .Y(G1218GAT_62_ngat) );
INVXL U_g2479 (.A(G1440GAT_334_gat), .Y(G1440GAT_334_ngat) );
INVXL U_g2480 (.A(G1170GAT_78_gat), .Y(G1170GAT_78_ngat) );
INVXL U_g2481 (.A(G1437GAT_335_gat), .Y(G1437GAT_335_ngat) );
INVXL U_g2482 (.A(G1122GAT_94_gat), .Y(G1122GAT_94_ngat) );
INVXL U_g2483 (.A(G1434GAT_336_gat), .Y(G1434GAT_336_ngat) );
INVXL U_g2484 (.A(G1074GAT_110_gat), .Y(G1074GAT_110_ngat) );
INVXL U_g2485 (.A(G1431GAT_337_gat), .Y(G1431GAT_337_ngat) );
INVXL U_g2486 (.A(G1026GAT_126_gat), .Y(G1026GAT_126_ngat) );
INVXL U_g2487 (.A(G1428GAT_338_gat), .Y(G1428GAT_338_ngat) );
INVXL U_g2488 (.A(G978GAT_142_gat), .Y(G978GAT_142_ngat) );
INVXL U_g2489 (.A(G1425GAT_339_gat), .Y(G1425GAT_339_ngat) );
INVXL U_g2490 (.A(G930GAT_158_gat), .Y(G930GAT_158_ngat) );
INVXL U_g2491 (.A(G1422GAT_340_gat), .Y(G1422GAT_340_ngat) );
INVXL U_g2492 (.A(G882GAT_174_gat), .Y(G882GAT_174_ngat) );
INVXL U_g2493 (.A(G1419GAT_341_gat), .Y(G1419GAT_341_ngat) );
INVXL U_g2494 (.A(G834GAT_190_gat), .Y(G834GAT_190_ngat) );
INVXL U_g2495 (.A(G1416GAT_342_gat), .Y(G1416GAT_342_ngat) );
INVXL U_g2496 (.A(G786GAT_206_gat), .Y(G786GAT_206_ngat) );
INVXL U_g2497 (.A(G1413GAT_343_gat), .Y(G1413GAT_343_ngat) );
INVXL U_g2498 (.A(G738GAT_222_gat), .Y(G738GAT_222_ngat) );
INVXL U_g2499 (.A(G1410GAT_344_gat), .Y(G1410GAT_344_ngat) );
INVXL U_g2500 (.A(G690GAT_238_gat), .Y(G690GAT_238_ngat) );
INVXL U_g2501 (.A(G1407GAT_345_gat), .Y(G1407GAT_345_ngat) );
INVXL U_g2502 (.A(G642GAT_254_gat), .Y(G642GAT_254_ngat) );
INVXL U_g2503 (.A(G1404GAT_346_gat), .Y(G1404GAT_346_ngat) );
INVXL U_g2504 (.A(G594GAT_270_gat), .Y(G594GAT_270_ngat) );
INVXL U_g2505 (.A(G1401GAT_347_gat), .Y(G1401GAT_347_ngat) );
INVXL U_g2506 (.A(G546GAT_286_gat), .Y(G546GAT_286_ngat) );
INVXL U_g2507 (.A(G1502GAT_348_gat), .Y(G1502GAT_348_ngat) );
INVXL U_g2508 (.A(G1498GAT_349_gat), .Y(G1498GAT_349_ngat) );
INVXL U_g2509 (.A(G1494GAT_350_gat), .Y(G1494GAT_350_ngat) );
INVXL U_g2510 (.A(G1490GAT_351_gat), .Y(G1490GAT_351_ngat) );
INVXL U_g2511 (.A(G1486GAT_352_gat), .Y(G1486GAT_352_ngat) );
INVXL U_g2512 (.A(G1482GAT_353_gat), .Y(G1482GAT_353_ngat) );
INVXL U_g2513 (.A(G1478GAT_354_gat), .Y(G1478GAT_354_ngat) );
INVXL U_g2514 (.A(G1474GAT_355_gat), .Y(G1474GAT_355_ngat) );
INVXL U_g2515 (.A(G1470GAT_356_gat), .Y(G1470GAT_356_ngat) );
INVXL U_g2516 (.A(G1466GAT_357_gat), .Y(G1466GAT_357_ngat) );
INVXL U_g2517 (.A(G1462GAT_358_gat), .Y(G1462GAT_358_ngat) );
INVXL U_g2518 (.A(G1458GAT_359_gat), .Y(G1458GAT_359_ngat) );
INVXL U_g2519 (.A(G1454GAT_360_gat), .Y(G1454GAT_360_ngat) );
INVXL U_g2520 (.A(G1450GAT_361_gat), .Y(G1450GAT_361_ngat) );
INVXL U_g2521 (.A(G1446GAT_362_gat), .Y(G1446GAT_362_ngat) );
INVXL U_g2522 (.A(G1266GAT_46_gat), .Y(G1266GAT_46_ngat) );
INVXL U_g2523 (.A(G1578GAT_363_gat), .Y(G1578GAT_363_ngat) );
INVXL U_g2524 (.A(G1576GAT_364_gat), .Y(G1576GAT_364_ngat) );
INVXL U_g2525 (.A(G1577GAT_365_gat), .Y(G1577GAT_365_ngat) );
INVXL U_g2526 (.A(G1571GAT_367_gat), .Y(G1571GAT_367_ngat) );
INVXL U_g2527 (.A(G1572GAT_368_gat), .Y(G1572GAT_368_ngat) );
INVXL U_g2528 (.A(G1566GAT_370_gat), .Y(G1566GAT_370_ngat) );
INVXL U_g2529 (.A(G1567GAT_371_gat), .Y(G1567GAT_371_ngat) );
INVXL U_g2530 (.A(G1561GAT_373_gat), .Y(G1561GAT_373_ngat) );
INVXL U_g2531 (.A(G1562GAT_374_gat), .Y(G1562GAT_374_ngat) );
INVXL U_g2532 (.A(G1556GAT_376_gat), .Y(G1556GAT_376_ngat) );
INVXL U_g2533 (.A(G1557GAT_377_gat), .Y(G1557GAT_377_ngat) );
INVXL U_g2534 (.A(G1551GAT_379_gat), .Y(G1551GAT_379_ngat) );
INVXL U_g2535 (.A(G1552GAT_380_gat), .Y(G1552GAT_380_ngat) );
INVXL U_g2536 (.A(G1546GAT_382_gat), .Y(G1546GAT_382_ngat) );
INVXL U_g2537 (.A(G1547GAT_383_gat), .Y(G1547GAT_383_ngat) );
INVXL U_g2538 (.A(G1541GAT_385_gat), .Y(G1541GAT_385_ngat) );
INVXL U_g2539 (.A(G1542GAT_386_gat), .Y(G1542GAT_386_ngat) );
INVXL U_g2540 (.A(G1536GAT_388_gat), .Y(G1536GAT_388_ngat) );
INVXL U_g2541 (.A(G1537GAT_389_gat), .Y(G1537GAT_389_ngat) );
INVXL U_g2542 (.A(G1531GAT_391_gat), .Y(G1531GAT_391_ngat) );
INVXL U_g2543 (.A(G1532GAT_392_gat), .Y(G1532GAT_392_ngat) );
INVXL U_g2544 (.A(G1526GAT_394_gat), .Y(G1526GAT_394_ngat) );
INVXL U_g2545 (.A(G1527GAT_395_gat), .Y(G1527GAT_395_ngat) );
INVXL U_g2546 (.A(G1521GAT_397_gat), .Y(G1521GAT_397_ngat) );
INVXL U_g2547 (.A(G1522GAT_398_gat), .Y(G1522GAT_398_ngat) );
INVXL U_g2548 (.A(G1516GAT_400_gat), .Y(G1516GAT_400_ngat) );
INVXL U_g2549 (.A(G1517GAT_401_gat), .Y(G1517GAT_401_ngat) );
INVXL U_g2550 (.A(G1511GAT_403_gat), .Y(G1511GAT_403_ngat) );
INVXL U_g2551 (.A(G1512GAT_404_gat), .Y(G1512GAT_404_ngat) );
INVXL U_g2552 (.A(G1506GAT_406_gat), .Y(G1506GAT_406_ngat) );
INVXL U_g2553 (.A(G1507GAT_407_gat), .Y(G1507GAT_407_ngat) );
INVXL U_g2554 (.A(G1624GAT_408_gat), .Y(G1624GAT_408_ngat) );
INVXL U_g2555 (.A(G1621GAT_409_gat), .Y(G1621GAT_409_ngat) );
INVXL U_g2556 (.A(G1573GAT_366_gat), .Y(G1573GAT_366_ngat) );
INVXL U_g2557 (.A(G1618GAT_410_gat), .Y(G1618GAT_410_ngat) );
INVXL U_g2558 (.A(G1568GAT_369_gat), .Y(G1568GAT_369_ngat) );
INVXL U_g2559 (.A(G1615GAT_411_gat), .Y(G1615GAT_411_ngat) );
INVXL U_g2560 (.A(G1563GAT_372_gat), .Y(G1563GAT_372_ngat) );
INVXL U_g2561 (.A(G1612GAT_412_gat), .Y(G1612GAT_412_ngat) );
INVXL U_g2562 (.A(G1558GAT_375_gat), .Y(G1558GAT_375_ngat) );
INVXL U_g2563 (.A(G1609GAT_413_gat), .Y(G1609GAT_413_ngat) );
INVXL U_g2564 (.A(G1553GAT_378_gat), .Y(G1553GAT_378_ngat) );
INVXL U_g2565 (.A(G1606GAT_414_gat), .Y(G1606GAT_414_ngat) );
INVXL U_g2566 (.A(G1548GAT_381_gat), .Y(G1548GAT_381_ngat) );
INVXL U_g2567 (.A(G1603GAT_415_gat), .Y(G1603GAT_415_ngat) );
INVXL U_g2568 (.A(G1543GAT_384_gat), .Y(G1543GAT_384_ngat) );
INVXL U_g2569 (.A(G1600GAT_416_gat), .Y(G1600GAT_416_ngat) );
INVXL U_g2570 (.A(G1538GAT_387_gat), .Y(G1538GAT_387_ngat) );
INVXL U_g2571 (.A(G1597GAT_417_gat), .Y(G1597GAT_417_ngat) );
INVXL U_g2572 (.A(G1533GAT_390_gat), .Y(G1533GAT_390_ngat) );
INVXL U_g2573 (.A(G1594GAT_418_gat), .Y(G1594GAT_418_ngat) );
INVXL U_g2574 (.A(G1528GAT_393_gat), .Y(G1528GAT_393_ngat) );
INVXL U_g2575 (.A(G1591GAT_419_gat), .Y(G1591GAT_419_ngat) );
INVXL U_g2576 (.A(G1523GAT_396_gat), .Y(G1523GAT_396_ngat) );
INVXL U_g2577 (.A(G1588GAT_420_gat), .Y(G1588GAT_420_ngat) );
INVXL U_g2578 (.A(G1518GAT_399_gat), .Y(G1518GAT_399_ngat) );
INVXL U_g2579 (.A(G1585GAT_421_gat), .Y(G1585GAT_421_ngat) );
INVXL U_g2580 (.A(G1513GAT_402_gat), .Y(G1513GAT_402_ngat) );
INVXL U_g2581 (.A(G1582GAT_422_gat), .Y(G1582GAT_422_ngat) );
INVXL U_g2582 (.A(G1508GAT_405_gat), .Y(G1508GAT_405_ngat) );
INVXL U_g2583 (.A(G1684GAT_424_gat), .Y(G1684GAT_424_ngat) );
INVXL U_g2584 (.A(G1685GAT_425_gat), .Y(G1685GAT_425_ngat) );
INVXL U_g2585 (.A(G1680GAT_426_gat), .Y(G1680GAT_426_ngat) );
INVXL U_g2586 (.A(G1676GAT_427_gat), .Y(G1676GAT_427_ngat) );
INVXL U_g2587 (.A(G1672GAT_428_gat), .Y(G1672GAT_428_ngat) );
INVXL U_g2588 (.A(G1668GAT_429_gat), .Y(G1668GAT_429_ngat) );
INVXL U_g2589 (.A(G1664GAT_430_gat), .Y(G1664GAT_430_ngat) );
INVXL U_g2590 (.A(G1660GAT_431_gat), .Y(G1660GAT_431_ngat) );
INVXL U_g2591 (.A(G1656GAT_432_gat), .Y(G1656GAT_432_ngat) );
INVXL U_g2592 (.A(G1652GAT_433_gat), .Y(G1652GAT_433_ngat) );
INVXL U_g2593 (.A(G1648GAT_434_gat), .Y(G1648GAT_434_ngat) );
INVXL U_g2594 (.A(G1644GAT_435_gat), .Y(G1644GAT_435_ngat) );
INVXL U_g2595 (.A(G1640GAT_436_gat), .Y(G1640GAT_436_ngat) );
INVXL U_g2596 (.A(G1636GAT_437_gat), .Y(G1636GAT_437_ngat) );
INVXL U_g2597 (.A(G1632GAT_438_gat), .Y(G1632GAT_438_ngat) );
INVXL U_g2598 (.A(G1628GAT_439_gat), .Y(G1628GAT_439_ngat) );
INVXL U_g2599 (.A(G1712GAT_441_gat), .Y(G1712GAT_441_ngat) );
INVXL U_g2600 (.A(G1713GAT_442_gat), .Y(G1713GAT_442_ngat) );
INVXL U_g2601 (.A(G1714GAT_440_gat), .Y(G1714GAT_440_ngat) );
INVXL U_g2602 (.A(G1221GAT_61_gat), .Y(G1221GAT_61_ngat) );
INVXL U_g2603 (.A(G1710GAT_443_gat), .Y(G1710GAT_443_ngat) );
INVXL U_g2604 (.A(G1711GAT_444_gat), .Y(G1711GAT_444_ngat) );
INVXL U_g2605 (.A(G1708GAT_445_gat), .Y(G1708GAT_445_ngat) );
INVXL U_g2606 (.A(G1709GAT_446_gat), .Y(G1709GAT_446_ngat) );
INVXL U_g2607 (.A(G1706GAT_447_gat), .Y(G1706GAT_447_ngat) );
INVXL U_g2608 (.A(G1707GAT_448_gat), .Y(G1707GAT_448_ngat) );
INVXL U_g2609 (.A(G1704GAT_449_gat), .Y(G1704GAT_449_ngat) );
INVXL U_g2610 (.A(G1705GAT_450_gat), .Y(G1705GAT_450_ngat) );
INVXL U_g2611 (.A(G1702GAT_451_gat), .Y(G1702GAT_451_ngat) );
INVXL U_g2612 (.A(G1703GAT_452_gat), .Y(G1703GAT_452_ngat) );
INVXL U_g2613 (.A(G1700GAT_453_gat), .Y(G1700GAT_453_ngat) );
INVXL U_g2614 (.A(G1701GAT_454_gat), .Y(G1701GAT_454_ngat) );
INVXL U_g2615 (.A(G1698GAT_455_gat), .Y(G1698GAT_455_ngat) );
INVXL U_g2616 (.A(G1699GAT_456_gat), .Y(G1699GAT_456_ngat) );
INVXL U_g2617 (.A(G1696GAT_457_gat), .Y(G1696GAT_457_ngat) );
INVXL U_g2618 (.A(G1697GAT_458_gat), .Y(G1697GAT_458_ngat) );
INVXL U_g2619 (.A(G1694GAT_459_gat), .Y(G1694GAT_459_ngat) );
INVXL U_g2620 (.A(G1695GAT_460_gat), .Y(G1695GAT_460_ngat) );
INVXL U_g2621 (.A(G1692GAT_461_gat), .Y(G1692GAT_461_ngat) );
INVXL U_g2622 (.A(G1693GAT_462_gat), .Y(G1693GAT_462_ngat) );
INVXL U_g2623 (.A(G1690GAT_463_gat), .Y(G1690GAT_463_ngat) );
INVXL U_g2624 (.A(G1691GAT_464_gat), .Y(G1691GAT_464_ngat) );
INVXL U_g2625 (.A(G1688GAT_465_gat), .Y(G1688GAT_465_ngat) );
INVXL U_g2626 (.A(G1689GAT_466_gat), .Y(G1689GAT_466_ngat) );
INVXL U_g2627 (.A(G1686GAT_467_gat), .Y(G1686GAT_467_ngat) );
INVXL U_g2628 (.A(G1687GAT_468_gat), .Y(G1687GAT_468_ngat) );
INVXL U_g2629 (.A(G1759GAT_470_gat), .Y(G1759GAT_470_ngat) );
INVXL U_g2630 (.A(G1756GAT_469_gat), .Y(G1756GAT_469_ngat) );
INVXL U_g2631 (.A(G1173GAT_77_gat), .Y(G1173GAT_77_ngat) );
INVXL U_g2632 (.A(G1753GAT_471_gat), .Y(G1753GAT_471_ngat) );
INVXL U_g2633 (.A(G1125GAT_93_gat), .Y(G1125GAT_93_ngat) );
INVXL U_g2634 (.A(G1750GAT_472_gat), .Y(G1750GAT_472_ngat) );
INVXL U_g2635 (.A(G1077GAT_109_gat), .Y(G1077GAT_109_ngat) );
INVXL U_g2636 (.A(G1747GAT_473_gat), .Y(G1747GAT_473_ngat) );
INVXL U_g2637 (.A(G1029GAT_125_gat), .Y(G1029GAT_125_ngat) );
INVXL U_g2638 (.A(G1744GAT_474_gat), .Y(G1744GAT_474_ngat) );
INVXL U_g2639 (.A(G981GAT_141_gat), .Y(G981GAT_141_ngat) );
INVXL U_g2640 (.A(G1741GAT_475_gat), .Y(G1741GAT_475_ngat) );
INVXL U_g2641 (.A(G933GAT_157_gat), .Y(G933GAT_157_ngat) );
INVXL U_g2642 (.A(G1738GAT_476_gat), .Y(G1738GAT_476_ngat) );
INVXL U_g2643 (.A(G885GAT_173_gat), .Y(G885GAT_173_ngat) );
INVXL U_g2644 (.A(G1735GAT_477_gat), .Y(G1735GAT_477_ngat) );
INVXL U_g2645 (.A(G837GAT_189_gat), .Y(G837GAT_189_ngat) );
INVXL U_g2646 (.A(G1732GAT_478_gat), .Y(G1732GAT_478_ngat) );
INVXL U_g2647 (.A(G789GAT_205_gat), .Y(G789GAT_205_ngat) );
INVXL U_g2648 (.A(G1729GAT_479_gat), .Y(G1729GAT_479_ngat) );
INVXL U_g2649 (.A(G741GAT_221_gat), .Y(G741GAT_221_ngat) );
INVXL U_g2650 (.A(G1726GAT_480_gat), .Y(G1726GAT_480_ngat) );
INVXL U_g2651 (.A(G693GAT_237_gat), .Y(G693GAT_237_ngat) );
INVXL U_g2652 (.A(G1723GAT_481_gat), .Y(G1723GAT_481_ngat) );
INVXL U_g2653 (.A(G645GAT_253_gat), .Y(G645GAT_253_ngat) );
INVXL U_g2654 (.A(G1720GAT_482_gat), .Y(G1720GAT_482_ngat) );
INVXL U_g2655 (.A(G597GAT_269_gat), .Y(G597GAT_269_ngat) );
INVXL U_g2656 (.A(G1717GAT_483_gat), .Y(G1717GAT_483_ngat) );
INVXL U_g2657 (.A(G549GAT_285_gat), .Y(G549GAT_285_ngat) );
INVXL U_g2658 (.A(G1269GAT_45_gat), .Y(G1269GAT_45_ngat) );
INVXL U_g2659 (.A(G1821GAT_484_gat), .Y(G1821GAT_484_ngat) );
INVXL U_g2660 (.A(G1819GAT_485_gat), .Y(G1819GAT_485_ngat) );
INVXL U_g2661 (.A(G1820GAT_486_gat), .Y(G1820GAT_486_ngat) );
INVXL U_g2662 (.A(G1815GAT_487_gat), .Y(G1815GAT_487_ngat) );
INVXL U_g2663 (.A(G1811GAT_488_gat), .Y(G1811GAT_488_ngat) );
INVXL U_g2664 (.A(G1807GAT_489_gat), .Y(G1807GAT_489_ngat) );
INVXL U_g2665 (.A(G1803GAT_490_gat), .Y(G1803GAT_490_ngat) );
INVXL U_g2666 (.A(G1799GAT_491_gat), .Y(G1799GAT_491_ngat) );
INVXL U_g2667 (.A(G1795GAT_492_gat), .Y(G1795GAT_492_ngat) );
INVXL U_g2668 (.A(G1791GAT_493_gat), .Y(G1791GAT_493_ngat) );
INVXL U_g2669 (.A(G1787GAT_494_gat), .Y(G1787GAT_494_ngat) );
INVXL U_g2670 (.A(G1783GAT_495_gat), .Y(G1783GAT_495_ngat) );
INVXL U_g2671 (.A(G1779GAT_496_gat), .Y(G1779GAT_496_ngat) );
INVXL U_g2672 (.A(G1775GAT_497_gat), .Y(G1775GAT_497_ngat) );
INVXL U_g2673 (.A(G1771GAT_498_gat), .Y(G1771GAT_498_ngat) );
INVXL U_g2674 (.A(G1767GAT_499_gat), .Y(G1767GAT_499_ngat) );
INVXL U_g2675 (.A(G1763GAT_500_gat), .Y(G1763GAT_500_ngat) );
INVXL U_g2676 (.A(G1897GAT_501_gat), .Y(G1897GAT_501_ngat) );
INVXL U_g2677 (.A(G1894GAT_502_gat), .Y(G1894GAT_502_ngat) );
INVXL U_g2678 (.A(G1891GAT_504_gat), .Y(G1891GAT_504_ngat) );
INVXL U_g2679 (.A(G1889GAT_503_gat), .Y(G1889GAT_503_ngat) );
INVXL U_g2680 (.A(G1890GAT_506_gat), .Y(G1890GAT_506_ngat) );
INVXL U_g2681 (.A(G1884GAT_505_gat), .Y(G1884GAT_505_ngat) );
INVXL U_g2682 (.A(G1885GAT_509_gat), .Y(G1885GAT_509_ngat) );
INVXL U_g2683 (.A(G1879GAT_508_gat), .Y(G1879GAT_508_ngat) );
INVXL U_g2684 (.A(G1880GAT_512_gat), .Y(G1880GAT_512_ngat) );
INVXL U_g2685 (.A(G1874GAT_511_gat), .Y(G1874GAT_511_ngat) );
INVXL U_g2686 (.A(G1875GAT_515_gat), .Y(G1875GAT_515_ngat) );
INVXL U_g2687 (.A(G1869GAT_514_gat), .Y(G1869GAT_514_ngat) );
INVXL U_g2688 (.A(G1870GAT_518_gat), .Y(G1870GAT_518_ngat) );
INVXL U_g2689 (.A(G1864GAT_517_gat), .Y(G1864GAT_517_ngat) );
INVXL U_g2690 (.A(G1865GAT_521_gat), .Y(G1865GAT_521_ngat) );
INVXL U_g2691 (.A(G1859GAT_520_gat), .Y(G1859GAT_520_ngat) );
INVXL U_g2692 (.A(G1860GAT_524_gat), .Y(G1860GAT_524_ngat) );
INVXL U_g2693 (.A(G1854GAT_523_gat), .Y(G1854GAT_523_ngat) );
INVXL U_g2694 (.A(G1855GAT_527_gat), .Y(G1855GAT_527_ngat) );
INVXL U_g2695 (.A(G1849GAT_526_gat), .Y(G1849GAT_526_ngat) );
INVXL U_g2696 (.A(G1850GAT_530_gat), .Y(G1850GAT_530_ngat) );
INVXL U_g2697 (.A(G1844GAT_529_gat), .Y(G1844GAT_529_ngat) );
INVXL U_g2698 (.A(G1845GAT_533_gat), .Y(G1845GAT_533_ngat) );
INVXL U_g2699 (.A(G1839GAT_532_gat), .Y(G1839GAT_532_ngat) );
INVXL U_g2700 (.A(G1840GAT_536_gat), .Y(G1840GAT_536_ngat) );
INVXL U_g2701 (.A(G1834GAT_535_gat), .Y(G1834GAT_535_ngat) );
INVXL U_g2702 (.A(G1835GAT_539_gat), .Y(G1835GAT_539_ngat) );
INVXL U_g2703 (.A(G1829GAT_538_gat), .Y(G1829GAT_538_ngat) );
INVXL U_g2704 (.A(G1830GAT_542_gat), .Y(G1830GAT_542_ngat) );
INVXL U_g2705 (.A(G1824GAT_541_gat), .Y(G1824GAT_541_ngat) );
INVXL U_g2706 (.A(G1825GAT_544_gat), .Y(G1825GAT_544_ngat) );
INVXL U_g2707 (.A(G1945GAT_545_gat), .Y(G1945GAT_545_ngat) );
INVXL U_g2708 (.A(G1946GAT_546_gat), .Y(G1946GAT_546_ngat) );
INVXL U_g2709 (.A(G1941GAT_547_gat), .Y(G1941GAT_547_ngat) );
INVXL U_g2710 (.A(G1938GAT_548_gat), .Y(G1938GAT_548_ngat) );
INVXL U_g2711 (.A(G1886GAT_507_gat), .Y(G1886GAT_507_ngat) );
INVXL U_g2712 (.A(G1935GAT_549_gat), .Y(G1935GAT_549_ngat) );
INVXL U_g2713 (.A(G1881GAT_510_gat), .Y(G1881GAT_510_ngat) );
INVXL U_g2714 (.A(G1932GAT_550_gat), .Y(G1932GAT_550_ngat) );
INVXL U_g2715 (.A(G1876GAT_513_gat), .Y(G1876GAT_513_ngat) );
INVXL U_g2716 (.A(G1929GAT_551_gat), .Y(G1929GAT_551_ngat) );
INVXL U_g2717 (.A(G1871GAT_516_gat), .Y(G1871GAT_516_ngat) );
INVXL U_g2718 (.A(G1926GAT_552_gat), .Y(G1926GAT_552_ngat) );
INVXL U_g2719 (.A(G1866GAT_519_gat), .Y(G1866GAT_519_ngat) );
INVXL U_g2720 (.A(G1923GAT_553_gat), .Y(G1923GAT_553_ngat) );
INVXL U_g2721 (.A(G1861GAT_522_gat), .Y(G1861GAT_522_ngat) );
INVXL U_g2722 (.A(G1920GAT_554_gat), .Y(G1920GAT_554_ngat) );
INVXL U_g2723 (.A(G1856GAT_525_gat), .Y(G1856GAT_525_ngat) );
INVXL U_g2724 (.A(G1917GAT_555_gat), .Y(G1917GAT_555_ngat) );
INVXL U_g2725 (.A(G1851GAT_528_gat), .Y(G1851GAT_528_ngat) );
INVXL U_g2726 (.A(G1914GAT_556_gat), .Y(G1914GAT_556_ngat) );
INVXL U_g2727 (.A(G1846GAT_531_gat), .Y(G1846GAT_531_ngat) );
INVXL U_g2728 (.A(G1911GAT_557_gat), .Y(G1911GAT_557_ngat) );
INVXL U_g2729 (.A(G1841GAT_534_gat), .Y(G1841GAT_534_ngat) );
INVXL U_g2730 (.A(G1908GAT_558_gat), .Y(G1908GAT_558_ngat) );
INVXL U_g2731 (.A(G1836GAT_537_gat), .Y(G1836GAT_537_ngat) );
INVXL U_g2732 (.A(G1905GAT_559_gat), .Y(G1905GAT_559_ngat) );
INVXL U_g2733 (.A(G1831GAT_540_gat), .Y(G1831GAT_540_ngat) );
INVXL U_g2734 (.A(G1902GAT_560_gat), .Y(G1902GAT_560_ngat) );
INVXL U_g2735 (.A(G1826GAT_543_gat), .Y(G1826GAT_543_ngat) );
INVXL U_g2736 (.A(G1999GAT_563_gat), .Y(G1999GAT_563_ngat) );
INVXL U_g2737 (.A(G2000GAT_564_gat), .Y(G2000GAT_564_ngat) );
INVXL U_g2738 (.A(G1995GAT_565_gat), .Y(G1995GAT_565_ngat) );
INVXL U_g2739 (.A(G2001GAT_562_gat), .Y(G2001GAT_562_ngat) );
INVXL U_g2740 (.A(G1224GAT_60_gat), .Y(G1224GAT_60_ngat) );
INVXL U_g2741 (.A(G1991GAT_566_gat), .Y(G1991GAT_566_ngat) );
INVXL U_g2742 (.A(G1987GAT_567_gat), .Y(G1987GAT_567_ngat) );
INVXL U_g2743 (.A(G1983GAT_568_gat), .Y(G1983GAT_568_ngat) );
INVXL U_g2744 (.A(G1979GAT_569_gat), .Y(G1979GAT_569_ngat) );
INVXL U_g2745 (.A(G1975GAT_570_gat), .Y(G1975GAT_570_ngat) );
INVXL U_g2746 (.A(G1971GAT_571_gat), .Y(G1971GAT_571_ngat) );
INVXL U_g2747 (.A(G1967GAT_572_gat), .Y(G1967GAT_572_ngat) );
INVXL U_g2748 (.A(G1963GAT_573_gat), .Y(G1963GAT_573_ngat) );
INVXL U_g2749 (.A(G1959GAT_574_gat), .Y(G1959GAT_574_ngat) );
INVXL U_g2750 (.A(G1955GAT_575_gat), .Y(G1955GAT_575_ngat) );
INVXL U_g2751 (.A(G1951GAT_576_gat), .Y(G1951GAT_576_ngat) );
INVXL U_g2752 (.A(G1947GAT_577_gat), .Y(G1947GAT_577_ngat) );
INVXL U_g2753 (.A(G2033GAT_580_gat), .Y(G2033GAT_580_ngat) );
INVXL U_g2754 (.A(G2028GAT_579_gat), .Y(G2028GAT_579_ngat) );
INVXL U_g2755 (.A(G2029GAT_582_gat), .Y(G2029GAT_582_ngat) );
INVXL U_g2756 (.A(G2026GAT_581_gat), .Y(G2026GAT_581_ngat) );
INVXL U_g2757 (.A(G2027GAT_584_gat), .Y(G2027GAT_584_ngat) );
INVXL U_g2758 (.A(G2030GAT_578_gat), .Y(G2030GAT_578_ngat) );
INVXL U_g2759 (.A(G1176GAT_76_gat), .Y(G1176GAT_76_ngat) );
INVXL U_g2760 (.A(G2024GAT_583_gat), .Y(G2024GAT_583_ngat) );
INVXL U_g2761 (.A(G2025GAT_586_gat), .Y(G2025GAT_586_ngat) );
INVXL U_g2762 (.A(G2022GAT_585_gat), .Y(G2022GAT_585_ngat) );
INVXL U_g2763 (.A(G2023GAT_588_gat), .Y(G2023GAT_588_ngat) );
INVXL U_g2764 (.A(G2020GAT_587_gat), .Y(G2020GAT_587_ngat) );
INVXL U_g2765 (.A(G2021GAT_590_gat), .Y(G2021GAT_590_ngat) );
INVXL U_g2766 (.A(G2018GAT_589_gat), .Y(G2018GAT_589_ngat) );
INVXL U_g2767 (.A(G2019GAT_592_gat), .Y(G2019GAT_592_ngat) );
INVXL U_g2768 (.A(G2016GAT_591_gat), .Y(G2016GAT_591_ngat) );
INVXL U_g2769 (.A(G2017GAT_594_gat), .Y(G2017GAT_594_ngat) );
INVXL U_g2770 (.A(G2014GAT_593_gat), .Y(G2014GAT_593_ngat) );
INVXL U_g2771 (.A(G2015GAT_596_gat), .Y(G2015GAT_596_ngat) );
INVXL U_g2772 (.A(G2012GAT_595_gat), .Y(G2012GAT_595_ngat) );
INVXL U_g2773 (.A(G2013GAT_598_gat), .Y(G2013GAT_598_ngat) );
INVXL U_g2774 (.A(G2010GAT_597_gat), .Y(G2010GAT_597_ngat) );
INVXL U_g2775 (.A(G2011GAT_600_gat), .Y(G2011GAT_600_ngat) );
INVXL U_g2776 (.A(G2008GAT_599_gat), .Y(G2008GAT_599_ngat) );
INVXL U_g2777 (.A(G2009GAT_602_gat), .Y(G2009GAT_602_ngat) );
INVXL U_g2778 (.A(G2006GAT_601_gat), .Y(G2006GAT_601_ngat) );
INVXL U_g2779 (.A(G2007GAT_604_gat), .Y(G2007GAT_604_ngat) );
INVXL U_g2780 (.A(G2004GAT_603_gat), .Y(G2004GAT_603_ngat) );
INVXL U_g2781 (.A(G2005GAT_605_gat), .Y(G2005GAT_605_ngat) );
INVXL U_g2782 (.A(G1272GAT_44_gat), .Y(G1272GAT_44_ngat) );
INVXL U_g2783 (.A(G2082GAT_606_gat), .Y(G2082GAT_606_ngat) );
INVXL U_g2784 (.A(G2080GAT_607_gat), .Y(G2080GAT_607_ngat) );
INVXL U_g2785 (.A(G2081GAT_609_gat), .Y(G2081GAT_609_ngat) );
INVXL U_g2786 (.A(G2076GAT_611_gat), .Y(G2076GAT_611_ngat) );
INVXL U_g2787 (.A(G2073GAT_608_gat), .Y(G2073GAT_608_ngat) );
INVXL U_g2788 (.A(G1128GAT_92_gat), .Y(G1128GAT_92_ngat) );
INVXL U_g2789 (.A(G2070GAT_610_gat), .Y(G2070GAT_610_ngat) );
INVXL U_g2790 (.A(G1080GAT_108_gat), .Y(G1080GAT_108_ngat) );
INVXL U_g2791 (.A(G2067GAT_612_gat), .Y(G2067GAT_612_ngat) );
INVXL U_g2792 (.A(G1032GAT_124_gat), .Y(G1032GAT_124_ngat) );
INVXL U_g2793 (.A(G2064GAT_613_gat), .Y(G2064GAT_613_ngat) );
INVXL U_g2794 (.A(G984GAT_140_gat), .Y(G984GAT_140_ngat) );
INVXL U_g2795 (.A(G2061GAT_614_gat), .Y(G2061GAT_614_ngat) );
INVXL U_g2796 (.A(G936GAT_156_gat), .Y(G936GAT_156_ngat) );
INVXL U_g2797 (.A(G2058GAT_615_gat), .Y(G2058GAT_615_ngat) );
INVXL U_g2798 (.A(G888GAT_172_gat), .Y(G888GAT_172_ngat) );
INVXL U_g2799 (.A(G2055GAT_616_gat), .Y(G2055GAT_616_ngat) );
INVXL U_g2800 (.A(G840GAT_188_gat), .Y(G840GAT_188_ngat) );
INVXL U_g2801 (.A(G2052GAT_617_gat), .Y(G2052GAT_617_ngat) );
INVXL U_g2802 (.A(G792GAT_204_gat), .Y(G792GAT_204_ngat) );
INVXL U_g2803 (.A(G2049GAT_618_gat), .Y(G2049GAT_618_ngat) );
INVXL U_g2804 (.A(G744GAT_220_gat), .Y(G744GAT_220_ngat) );
INVXL U_g2805 (.A(G2046GAT_619_gat), .Y(G2046GAT_619_ngat) );
INVXL U_g2806 (.A(G696GAT_236_gat), .Y(G696GAT_236_ngat) );
INVXL U_g2807 (.A(G2043GAT_620_gat), .Y(G2043GAT_620_ngat) );
INVXL U_g2808 (.A(G648GAT_252_gat), .Y(G648GAT_252_ngat) );
INVXL U_g2809 (.A(G2040GAT_621_gat), .Y(G2040GAT_621_ngat) );
INVXL U_g2810 (.A(G600GAT_268_gat), .Y(G600GAT_268_ngat) );
INVXL U_g2811 (.A(G2037GAT_622_gat), .Y(G2037GAT_622_ngat) );
INVXL U_g2812 (.A(G552GAT_284_gat), .Y(G552GAT_284_ngat) );
INVXL U_g2813 (.A(G2145GAT_623_gat), .Y(G2145GAT_623_ngat) );
INVXL U_g2814 (.A(G2142GAT_624_gat), .Y(G2142GAT_624_ngat) );
INVXL U_g2815 (.A(G2139GAT_625_gat), .Y(G2139GAT_625_ngat) );
INVXL U_g2816 (.A(G2137GAT_626_gat), .Y(G2137GAT_626_ngat) );
INVXL U_g2817 (.A(G2138GAT_627_gat), .Y(G2138GAT_627_ngat) );
INVXL U_g2818 (.A(G2133GAT_628_gat), .Y(G2133GAT_628_ngat) );
INVXL U_g2819 (.A(G2129GAT_629_gat), .Y(G2129GAT_629_ngat) );
INVXL U_g2820 (.A(G2125GAT_630_gat), .Y(G2125GAT_630_ngat) );
INVXL U_g2821 (.A(G2121GAT_631_gat), .Y(G2121GAT_631_ngat) );
INVXL U_g2822 (.A(G2117GAT_632_gat), .Y(G2117GAT_632_ngat) );
INVXL U_g2823 (.A(G2113GAT_633_gat), .Y(G2113GAT_633_ngat) );
INVXL U_g2824 (.A(G2109GAT_634_gat), .Y(G2109GAT_634_ngat) );
INVXL U_g2825 (.A(G2105GAT_635_gat), .Y(G2105GAT_635_ngat) );
INVXL U_g2826 (.A(G2101GAT_636_gat), .Y(G2101GAT_636_ngat) );
INVXL U_g2827 (.A(G2097GAT_637_gat), .Y(G2097GAT_637_ngat) );
INVXL U_g2828 (.A(G2093GAT_638_gat), .Y(G2093GAT_638_ngat) );
INVXL U_g2829 (.A(G2089GAT_639_gat), .Y(G2089GAT_639_ngat) );
INVXL U_g2830 (.A(G2085GAT_640_gat), .Y(G2085GAT_640_ngat) );
INVXL U_g2831 (.A(G2221GAT_641_gat), .Y(G2221GAT_641_ngat) );
INVXL U_g2832 (.A(G2222GAT_642_gat), .Y(G2222GAT_642_ngat) );
INVXL U_g2833 (.A(G2217GAT_643_gat), .Y(G2217GAT_643_ngat) );
INVXL U_g2834 (.A(G2214GAT_644_gat), .Y(G2214GAT_644_ngat) );
INVXL U_g2835 (.A(G2211GAT_647_gat), .Y(G2211GAT_647_ngat) );
INVXL U_g2836 (.A(G2209GAT_645_gat), .Y(G2209GAT_645_ngat) );
INVXL U_g2837 (.A(G2210GAT_649_gat), .Y(G2210GAT_649_ngat) );
INVXL U_g2838 (.A(G2204GAT_646_gat), .Y(G2204GAT_646_ngat) );
INVXL U_g2839 (.A(G2205GAT_652_gat), .Y(G2205GAT_652_ngat) );
INVXL U_g2840 (.A(G2199GAT_648_gat), .Y(G2199GAT_648_ngat) );
INVXL U_g2841 (.A(G2200GAT_655_gat), .Y(G2200GAT_655_ngat) );
INVXL U_g2842 (.A(G2194GAT_651_gat), .Y(G2194GAT_651_ngat) );
INVXL U_g2843 (.A(G2195GAT_658_gat), .Y(G2195GAT_658_ngat) );
INVXL U_g2844 (.A(G2189GAT_654_gat), .Y(G2189GAT_654_ngat) );
INVXL U_g2845 (.A(G2190GAT_661_gat), .Y(G2190GAT_661_ngat) );
INVXL U_g2846 (.A(G2184GAT_657_gat), .Y(G2184GAT_657_ngat) );
INVXL U_g2847 (.A(G2185GAT_664_gat), .Y(G2185GAT_664_ngat) );
INVXL U_g2848 (.A(G2179GAT_660_gat), .Y(G2179GAT_660_ngat) );
INVXL U_g2849 (.A(G2180GAT_667_gat), .Y(G2180GAT_667_ngat) );
INVXL U_g2850 (.A(G2174GAT_663_gat), .Y(G2174GAT_663_ngat) );
INVXL U_g2851 (.A(G2175GAT_670_gat), .Y(G2175GAT_670_ngat) );
INVXL U_g2852 (.A(G2169GAT_666_gat), .Y(G2169GAT_666_ngat) );
INVXL U_g2853 (.A(G2170GAT_673_gat), .Y(G2170GAT_673_ngat) );
INVXL U_g2854 (.A(G2164GAT_669_gat), .Y(G2164GAT_669_ngat) );
INVXL U_g2855 (.A(G2165GAT_676_gat), .Y(G2165GAT_676_ngat) );
INVXL U_g2856 (.A(G2159GAT_672_gat), .Y(G2159GAT_672_ngat) );
INVXL U_g2857 (.A(G2160GAT_679_gat), .Y(G2160GAT_679_ngat) );
INVXL U_g2858 (.A(G2154GAT_675_gat), .Y(G2154GAT_675_ngat) );
INVXL U_g2859 (.A(G2155GAT_681_gat), .Y(G2155GAT_681_ngat) );
INVXL U_g2860 (.A(G2149GAT_678_gat), .Y(G2149GAT_678_ngat) );
INVXL U_g2861 (.A(G2150GAT_683_gat), .Y(G2150GAT_683_ngat) );
INVXL U_g2862 (.A(G2264GAT_685_gat), .Y(G2264GAT_685_ngat) );
INVXL U_g2863 (.A(G2265GAT_686_gat), .Y(G2265GAT_686_ngat) );
INVXL U_g2864 (.A(G2260GAT_687_gat), .Y(G2260GAT_687_ngat) );
INVXL U_g2865 (.A(G2266GAT_684_gat), .Y(G2266GAT_684_ngat) );
INVXL U_g2866 (.A(G1227GAT_59_gat), .Y(G1227GAT_59_ngat) );
INVXL U_g2867 (.A(G2257GAT_688_gat), .Y(G2257GAT_688_ngat) );
INVXL U_g2868 (.A(G2206GAT_650_gat), .Y(G2206GAT_650_ngat) );
INVXL U_g2869 (.A(G2254GAT_689_gat), .Y(G2254GAT_689_ngat) );
INVXL U_g2870 (.A(G2201GAT_653_gat), .Y(G2201GAT_653_ngat) );
INVXL U_g2871 (.A(G2251GAT_690_gat), .Y(G2251GAT_690_ngat) );
INVXL U_g2872 (.A(G2196GAT_656_gat), .Y(G2196GAT_656_ngat) );
INVXL U_g2873 (.A(G2248GAT_691_gat), .Y(G2248GAT_691_ngat) );
INVXL U_g2874 (.A(G2191GAT_659_gat), .Y(G2191GAT_659_ngat) );
INVXL U_g2875 (.A(G2245GAT_692_gat), .Y(G2245GAT_692_ngat) );
INVXL U_g2876 (.A(G2186GAT_662_gat), .Y(G2186GAT_662_ngat) );
INVXL U_g2877 (.A(G2242GAT_693_gat), .Y(G2242GAT_693_ngat) );
INVXL U_g2878 (.A(G2181GAT_665_gat), .Y(G2181GAT_665_ngat) );
INVXL U_g2879 (.A(G2239GAT_694_gat), .Y(G2239GAT_694_ngat) );
INVXL U_g2880 (.A(G2176GAT_668_gat), .Y(G2176GAT_668_ngat) );
INVXL U_g2881 (.A(G2236GAT_695_gat), .Y(G2236GAT_695_ngat) );
INVXL U_g2882 (.A(G2171GAT_671_gat), .Y(G2171GAT_671_ngat) );
INVXL U_g2883 (.A(G2233GAT_696_gat), .Y(G2233GAT_696_ngat) );
INVXL U_g2884 (.A(G2166GAT_674_gat), .Y(G2166GAT_674_ngat) );
INVXL U_g2885 (.A(G2230GAT_697_gat), .Y(G2230GAT_697_ngat) );
INVXL U_g2886 (.A(G2161GAT_677_gat), .Y(G2161GAT_677_ngat) );
INVXL U_g2887 (.A(G2227GAT_698_gat), .Y(G2227GAT_698_ngat) );
INVXL U_g2888 (.A(G2156GAT_680_gat), .Y(G2156GAT_680_ngat) );
INVXL U_g2889 (.A(G2224GAT_699_gat), .Y(G2224GAT_699_ngat) );
INVXL U_g2890 (.A(G2151GAT_682_gat), .Y(G2151GAT_682_ngat) );
INVXL U_g2891 (.A(G2322GAT_703_gat), .Y(G2322GAT_703_ngat) );
INVXL U_g2892 (.A(G2317GAT_702_gat), .Y(G2317GAT_702_ngat) );
INVXL U_g2893 (.A(G2318GAT_704_gat), .Y(G2318GAT_704_ngat) );
INVXL U_g2894 (.A(G2313GAT_705_gat), .Y(G2313GAT_705_ngat) );
INVXL U_g2895 (.A(G2309GAT_706_gat), .Y(G2309GAT_706_ngat) );
INVXL U_g2896 (.A(G2319GAT_701_gat), .Y(G2319GAT_701_ngat) );
INVXL U_g2897 (.A(G1179GAT_75_gat), .Y(G1179GAT_75_ngat) );
INVXL U_g2898 (.A(G2305GAT_707_gat), .Y(G2305GAT_707_ngat) );
INVXL U_g2899 (.A(G2301GAT_708_gat), .Y(G2301GAT_708_ngat) );
INVXL U_g2900 (.A(G2297GAT_709_gat), .Y(G2297GAT_709_ngat) );
INVXL U_g2901 (.A(G2293GAT_710_gat), .Y(G2293GAT_710_ngat) );
INVXL U_g2902 (.A(G2289GAT_711_gat), .Y(G2289GAT_711_ngat) );
INVXL U_g2903 (.A(G2285GAT_712_gat), .Y(G2285GAT_712_ngat) );
INVXL U_g2904 (.A(G2281GAT_713_gat), .Y(G2281GAT_713_ngat) );
INVXL U_g2905 (.A(G2277GAT_714_gat), .Y(G2277GAT_714_ngat) );
INVXL U_g2906 (.A(G2273GAT_715_gat), .Y(G2273GAT_715_ngat) );
INVXL U_g2907 (.A(G2269GAT_716_gat), .Y(G2269GAT_716_ngat) );
INVXL U_g2908 (.A(G1275GAT_43_gat), .Y(G1275GAT_43_ngat) );
INVXL U_g2909 (.A(G2359GAT_717_gat), .Y(G2359GAT_717_ngat) );
INVXL U_g2910 (.A(G2357GAT_718_gat), .Y(G2357GAT_718_ngat) );
INVXL U_g2911 (.A(G2358GAT_721_gat), .Y(G2358GAT_721_ngat) );
INVXL U_g2912 (.A(G2353GAT_723_gat), .Y(G2353GAT_723_ngat) );
INVXL U_g2913 (.A(G2348GAT_720_gat), .Y(G2348GAT_720_ngat) );
INVXL U_g2914 (.A(G2349GAT_725_gat), .Y(G2349GAT_725_ngat) );
INVXL U_g2915 (.A(G2346GAT_722_gat), .Y(G2346GAT_722_ngat) );
INVXL U_g2916 (.A(G2347GAT_727_gat), .Y(G2347GAT_727_ngat) );
INVXL U_g2917 (.A(G2344GAT_724_gat), .Y(G2344GAT_724_ngat) );
INVXL U_g2918 (.A(G2345GAT_729_gat), .Y(G2345GAT_729_ngat) );
INVXL U_g2919 (.A(G2350GAT_719_gat), .Y(G2350GAT_719_ngat) );
INVXL U_g2920 (.A(G1131GAT_91_gat), .Y(G1131GAT_91_ngat) );
INVXL U_g2921 (.A(G2342GAT_726_gat), .Y(G2342GAT_726_ngat) );
INVXL U_g2922 (.A(G2343GAT_731_gat), .Y(G2343GAT_731_ngat) );
INVXL U_g2923 (.A(G2340GAT_728_gat), .Y(G2340GAT_728_ngat) );
INVXL U_g2924 (.A(G2341GAT_733_gat), .Y(G2341GAT_733_ngat) );
INVXL U_g2925 (.A(G2338GAT_730_gat), .Y(G2338GAT_730_ngat) );
INVXL U_g2926 (.A(G2339GAT_735_gat), .Y(G2339GAT_735_ngat) );
INVXL U_g2927 (.A(G2336GAT_732_gat), .Y(G2336GAT_732_ngat) );
INVXL U_g2928 (.A(G2337GAT_737_gat), .Y(G2337GAT_737_ngat) );
INVXL U_g2929 (.A(G2334GAT_734_gat), .Y(G2334GAT_734_ngat) );
INVXL U_g2930 (.A(G2335GAT_739_gat), .Y(G2335GAT_739_ngat) );
INVXL U_g2931 (.A(G2332GAT_736_gat), .Y(G2332GAT_736_ngat) );
INVXL U_g2932 (.A(G2333GAT_741_gat), .Y(G2333GAT_741_ngat) );
INVXL U_g2933 (.A(G2330GAT_738_gat), .Y(G2330GAT_738_ngat) );
INVXL U_g2934 (.A(G2331GAT_743_gat), .Y(G2331GAT_743_ngat) );
INVXL U_g2935 (.A(G2328GAT_740_gat), .Y(G2328GAT_740_ngat) );
INVXL U_g2936 (.A(G2329GAT_744_gat), .Y(G2329GAT_744_ngat) );
INVXL U_g2937 (.A(G2326GAT_742_gat), .Y(G2326GAT_742_ngat) );
INVXL U_g2938 (.A(G2327GAT_745_gat), .Y(G2327GAT_745_ngat) );
INVXL U_g2939 (.A(G2410GAT_746_gat), .Y(G2410GAT_746_ngat) );
INVXL U_g2940 (.A(G2407GAT_747_gat), .Y(G2407GAT_747_ngat) );
INVXL U_g2941 (.A(G2404GAT_748_gat), .Y(G2404GAT_748_ngat) );
INVXL U_g2942 (.A(G2402GAT_749_gat), .Y(G2402GAT_749_ngat) );
INVXL U_g2943 (.A(G2403GAT_752_gat), .Y(G2403GAT_752_ngat) );
INVXL U_g2944 (.A(G2398GAT_754_gat), .Y(G2398GAT_754_ngat) );
INVXL U_g2945 (.A(G2395GAT_750_gat), .Y(G2395GAT_750_ngat) );
INVXL U_g2946 (.A(G1083GAT_107_gat), .Y(G1083GAT_107_ngat) );
INVXL U_g2947 (.A(G2392GAT_751_gat), .Y(G2392GAT_751_ngat) );
INVXL U_g2948 (.A(G1035GAT_123_gat), .Y(G1035GAT_123_ngat) );
INVXL U_g2949 (.A(G2389GAT_753_gat), .Y(G2389GAT_753_ngat) );
INVXL U_g2950 (.A(G987GAT_139_gat), .Y(G987GAT_139_ngat) );
INVXL U_g2951 (.A(G2386GAT_755_gat), .Y(G2386GAT_755_ngat) );
INVXL U_g2952 (.A(G939GAT_155_gat), .Y(G939GAT_155_ngat) );
INVXL U_g2953 (.A(G2383GAT_756_gat), .Y(G2383GAT_756_ngat) );
INVXL U_g2954 (.A(G891GAT_171_gat), .Y(G891GAT_171_ngat) );
INVXL U_g2955 (.A(G2380GAT_757_gat), .Y(G2380GAT_757_ngat) );
INVXL U_g2956 (.A(G843GAT_187_gat), .Y(G843GAT_187_ngat) );
INVXL U_g2957 (.A(G2377GAT_758_gat), .Y(G2377GAT_758_ngat) );
INVXL U_g2958 (.A(G795GAT_203_gat), .Y(G795GAT_203_ngat) );
INVXL U_g2959 (.A(G2374GAT_759_gat), .Y(G2374GAT_759_ngat) );
INVXL U_g2960 (.A(G747GAT_219_gat), .Y(G747GAT_219_ngat) );
INVXL U_g2961 (.A(G2371GAT_760_gat), .Y(G2371GAT_760_ngat) );
INVXL U_g2962 (.A(G699GAT_235_gat), .Y(G699GAT_235_ngat) );
INVXL U_g2963 (.A(G2368GAT_761_gat), .Y(G2368GAT_761_ngat) );
INVXL U_g2964 (.A(G651GAT_251_gat), .Y(G651GAT_251_ngat) );
INVXL U_g2965 (.A(G2365GAT_762_gat), .Y(G2365GAT_762_ngat) );
INVXL U_g2966 (.A(G603GAT_267_gat), .Y(G603GAT_267_ngat) );
INVXL U_g2967 (.A(G2362GAT_763_gat), .Y(G2362GAT_763_ngat) );
INVXL U_g2968 (.A(G555GAT_283_gat), .Y(G555GAT_283_ngat) );
INVXL U_g2969 (.A(G2474GAT_764_gat), .Y(G2474GAT_764_ngat) );
INVXL U_g2970 (.A(G2475GAT_765_gat), .Y(G2475GAT_765_ngat) );
INVXL U_g2971 (.A(G2470GAT_766_gat), .Y(G2470GAT_766_ngat) );
INVXL U_g2972 (.A(G2467GAT_767_gat), .Y(G2467GAT_767_ngat) );
INVXL U_g2973 (.A(G2464GAT_768_gat), .Y(G2464GAT_768_ngat) );
INVXL U_g2974 (.A(G2462GAT_769_gat), .Y(G2462GAT_769_ngat) );
INVXL U_g2975 (.A(G2463GAT_770_gat), .Y(G2463GAT_770_ngat) );
INVXL U_g2976 (.A(G2458GAT_771_gat), .Y(G2458GAT_771_ngat) );
INVXL U_g2977 (.A(G2454GAT_772_gat), .Y(G2454GAT_772_ngat) );
INVXL U_g2978 (.A(G2450GAT_773_gat), .Y(G2450GAT_773_ngat) );
INVXL U_g2979 (.A(G2446GAT_774_gat), .Y(G2446GAT_774_ngat) );
INVXL U_g2980 (.A(G2442GAT_775_gat), .Y(G2442GAT_775_ngat) );
INVXL U_g2981 (.A(G2438GAT_776_gat), .Y(G2438GAT_776_ngat) );
INVXL U_g2982 (.A(G2434GAT_777_gat), .Y(G2434GAT_777_ngat) );
INVXL U_g2983 (.A(G2430GAT_778_gat), .Y(G2430GAT_778_ngat) );
INVXL U_g2984 (.A(G2426GAT_779_gat), .Y(G2426GAT_779_ngat) );
INVXL U_g2985 (.A(G2422GAT_780_gat), .Y(G2422GAT_780_ngat) );
INVXL U_g2986 (.A(G2418GAT_781_gat), .Y(G2418GAT_781_ngat) );
INVXL U_g2987 (.A(G2414GAT_782_gat), .Y(G2414GAT_782_ngat) );
INVXL U_g2988 (.A(G2543GAT_784_gat), .Y(G2543GAT_784_ngat) );
INVXL U_g2989 (.A(G2544GAT_785_gat), .Y(G2544GAT_785_ngat) );
INVXL U_g2990 (.A(G2539GAT_786_gat), .Y(G2539GAT_786_ngat) );
INVXL U_g2991 (.A(G2536GAT_787_gat), .Y(G2536GAT_787_ngat) );
INVXL U_g2992 (.A(G2533GAT_791_gat), .Y(G2533GAT_791_ngat) );
INVXL U_g2993 (.A(G2531GAT_788_gat), .Y(G2531GAT_788_ngat) );
INVXL U_g2994 (.A(G2532GAT_793_gat), .Y(G2532GAT_793_ngat) );
INVXL U_g2995 (.A(G2545GAT_783_gat), .Y(G2545GAT_783_ngat) );
INVXL U_g2996 (.A(G1230GAT_58_gat), .Y(G1230GAT_58_ngat) );
INVXL U_g2997 (.A(G2526GAT_789_gat), .Y(G2526GAT_789_ngat) );
INVXL U_g2998 (.A(G2527GAT_796_gat), .Y(G2527GAT_796_ngat) );
INVXL U_g2999 (.A(G2521GAT_790_gat), .Y(G2521GAT_790_ngat) );
INVXL U_g3000 (.A(G2522GAT_799_gat), .Y(G2522GAT_799_ngat) );
INVXL U_g3001 (.A(G2516GAT_792_gat), .Y(G2516GAT_792_ngat) );
INVXL U_g3002 (.A(G2517GAT_802_gat), .Y(G2517GAT_802_ngat) );
INVXL U_g3003 (.A(G2511GAT_795_gat), .Y(G2511GAT_795_ngat) );
INVXL U_g3004 (.A(G2512GAT_805_gat), .Y(G2512GAT_805_ngat) );
INVXL U_g3005 (.A(G2506GAT_798_gat), .Y(G2506GAT_798_ngat) );
INVXL U_g3006 (.A(G2507GAT_808_gat), .Y(G2507GAT_808_ngat) );
INVXL U_g3007 (.A(G2501GAT_801_gat), .Y(G2501GAT_801_ngat) );
INVXL U_g3008 (.A(G2502GAT_811_gat), .Y(G2502GAT_811_ngat) );
INVXL U_g3009 (.A(G2496GAT_804_gat), .Y(G2496GAT_804_ngat) );
INVXL U_g3010 (.A(G2497GAT_814_gat), .Y(G2497GAT_814_ngat) );
INVXL U_g3011 (.A(G2491GAT_807_gat), .Y(G2491GAT_807_ngat) );
INVXL U_g3012 (.A(G2492GAT_817_gat), .Y(G2492GAT_817_ngat) );
INVXL U_g3013 (.A(G2486GAT_810_gat), .Y(G2486GAT_810_ngat) );
INVXL U_g3014 (.A(G2487GAT_819_gat), .Y(G2487GAT_819_ngat) );
INVXL U_g3015 (.A(G2481GAT_813_gat), .Y(G2481GAT_813_ngat) );
INVXL U_g3016 (.A(G2482GAT_821_gat), .Y(G2482GAT_821_ngat) );
INVXL U_g3017 (.A(G2476GAT_816_gat), .Y(G2476GAT_816_ngat) );
INVXL U_g3018 (.A(G2477GAT_823_gat), .Y(G2477GAT_823_ngat) );
INVXL U_g3019 (.A(G2591GAT_829_gat), .Y(G2591GAT_829_ngat) );
INVXL U_g3020 (.A(G2586GAT_825_gat), .Y(G2586GAT_825_ngat) );
INVXL U_g3021 (.A(G2587GAT_826_gat), .Y(G2587GAT_826_ngat) );
INVXL U_g3022 (.A(G2582GAT_827_gat), .Y(G2582GAT_827_ngat) );
INVXL U_g3023 (.A(G2588GAT_824_gat), .Y(G2588GAT_824_ngat) );
INVXL U_g3024 (.A(G1182GAT_74_gat), .Y(G1182GAT_74_ngat) );
INVXL U_g3025 (.A(G2579GAT_828_gat), .Y(G2579GAT_828_ngat) );
INVXL U_g3026 (.A(G2528GAT_794_gat), .Y(G2528GAT_794_ngat) );
INVXL U_g3027 (.A(G2576GAT_830_gat), .Y(G2576GAT_830_ngat) );
INVXL U_g3028 (.A(G2523GAT_797_gat), .Y(G2523GAT_797_ngat) );
INVXL U_g3029 (.A(G2573GAT_831_gat), .Y(G2573GAT_831_ngat) );
INVXL U_g3030 (.A(G2518GAT_800_gat), .Y(G2518GAT_800_ngat) );
INVXL U_g3031 (.A(G2570GAT_832_gat), .Y(G2570GAT_832_ngat) );
INVXL U_g3032 (.A(G2513GAT_803_gat), .Y(G2513GAT_803_ngat) );
INVXL U_g3033 (.A(G2567GAT_833_gat), .Y(G2567GAT_833_ngat) );
INVXL U_g3034 (.A(G2508GAT_806_gat), .Y(G2508GAT_806_ngat) );
INVXL U_g3035 (.A(G2564GAT_834_gat), .Y(G2564GAT_834_ngat) );
INVXL U_g3036 (.A(G2503GAT_809_gat), .Y(G2503GAT_809_ngat) );
INVXL U_g3037 (.A(G2561GAT_835_gat), .Y(G2561GAT_835_ngat) );
INVXL U_g3038 (.A(G2498GAT_812_gat), .Y(G2498GAT_812_ngat) );
INVXL U_g3039 (.A(G2558GAT_836_gat), .Y(G2558GAT_836_ngat) );
INVXL U_g3040 (.A(G2493GAT_815_gat), .Y(G2493GAT_815_ngat) );
INVXL U_g3041 (.A(G2555GAT_837_gat), .Y(G2555GAT_837_ngat) );
INVXL U_g3042 (.A(G2488GAT_818_gat), .Y(G2488GAT_818_ngat) );
INVXL U_g3043 (.A(G2552GAT_838_gat), .Y(G2552GAT_838_ngat) );
INVXL U_g3044 (.A(G2483GAT_820_gat), .Y(G2483GAT_820_ngat) );
INVXL U_g3045 (.A(G2549GAT_839_gat), .Y(G2549GAT_839_ngat) );
INVXL U_g3046 (.A(G2478GAT_822_gat), .Y(G2478GAT_822_ngat) );
INVXL U_g3047 (.A(G1278GAT_42_gat), .Y(G1278GAT_42_ngat) );
INVXL U_g3048 (.A(G2650GAT_841_gat), .Y(G2650GAT_841_ngat) );
INVXL U_g3049 (.A(G2648GAT_842_gat), .Y(G2648GAT_842_ngat) );
INVXL U_g3050 (.A(G2649GAT_845_gat), .Y(G2649GAT_845_ngat) );
INVXL U_g3051 (.A(G2644GAT_846_gat), .Y(G2644GAT_846_ngat) );
INVXL U_g3052 (.A(G2639GAT_844_gat), .Y(G2639GAT_844_ngat) );
INVXL U_g3053 (.A(G2640GAT_847_gat), .Y(G2640GAT_847_ngat) );
INVXL U_g3054 (.A(G2635GAT_848_gat), .Y(G2635GAT_848_ngat) );
INVXL U_g3055 (.A(G2631GAT_849_gat), .Y(G2631GAT_849_ngat) );
INVXL U_g3056 (.A(G2627GAT_850_gat), .Y(G2627GAT_850_ngat) );
INVXL U_g3057 (.A(G2641GAT_843_gat), .Y(G2641GAT_843_ngat) );
INVXL U_g3058 (.A(G1134GAT_90_gat), .Y(G1134GAT_90_ngat) );
INVXL U_g3059 (.A(G2623GAT_851_gat), .Y(G2623GAT_851_ngat) );
INVXL U_g3060 (.A(G2619GAT_852_gat), .Y(G2619GAT_852_ngat) );
INVXL U_g3061 (.A(G2615GAT_853_gat), .Y(G2615GAT_853_ngat) );
INVXL U_g3062 (.A(G2611GAT_854_gat), .Y(G2611GAT_854_ngat) );
INVXL U_g3063 (.A(G2607GAT_855_gat), .Y(G2607GAT_855_ngat) );
INVXL U_g3064 (.A(G2603GAT_856_gat), .Y(G2603GAT_856_ngat) );
INVXL U_g3065 (.A(G2599GAT_857_gat), .Y(G2599GAT_857_ngat) );
INVXL U_g3066 (.A(G2595GAT_858_gat), .Y(G2595GAT_858_ngat) );
INVXL U_g3067 (.A(G2690GAT_859_gat), .Y(G2690GAT_859_ngat) );
INVXL U_g3068 (.A(G2687GAT_860_gat), .Y(G2687GAT_860_ngat) );
INVXL U_g3069 (.A(G2684GAT_861_gat), .Y(G2684GAT_861_ngat) );
INVXL U_g3070 (.A(G2682GAT_862_gat), .Y(G2682GAT_862_ngat) );
INVXL U_g3071 (.A(G2683GAT_866_gat), .Y(G2683GAT_866_ngat) );
INVXL U_g3072 (.A(G2678GAT_868_gat), .Y(G2678GAT_868_ngat) );
INVXL U_g3073 (.A(G2673GAT_864_gat), .Y(G2673GAT_864_ngat) );
INVXL U_g3074 (.A(G2674GAT_870_gat), .Y(G2674GAT_870_ngat) );
INVXL U_g3075 (.A(G2671GAT_865_gat), .Y(G2671GAT_865_ngat) );
INVXL U_g3076 (.A(G2672GAT_872_gat), .Y(G2672GAT_872_ngat) );
INVXL U_g3077 (.A(G2669GAT_867_gat), .Y(G2669GAT_867_ngat) );
INVXL U_g3078 (.A(G2670GAT_874_gat), .Y(G2670GAT_874_ngat) );
INVXL U_g3079 (.A(G2667GAT_869_gat), .Y(G2667GAT_869_ngat) );
INVXL U_g3080 (.A(G2668GAT_876_gat), .Y(G2668GAT_876_ngat) );
INVXL U_g3081 (.A(G2675GAT_863_gat), .Y(G2675GAT_863_ngat) );
INVXL U_g3082 (.A(G1086GAT_106_gat), .Y(G1086GAT_106_ngat) );
INVXL U_g3083 (.A(G2665GAT_871_gat), .Y(G2665GAT_871_ngat) );
INVXL U_g3084 (.A(G2666GAT_878_gat), .Y(G2666GAT_878_ngat) );
INVXL U_g3085 (.A(G2663GAT_873_gat), .Y(G2663GAT_873_ngat) );
INVXL U_g3086 (.A(G2664GAT_880_gat), .Y(G2664GAT_880_ngat) );
INVXL U_g3087 (.A(G2661GAT_875_gat), .Y(G2661GAT_875_ngat) );
INVXL U_g3088 (.A(G2662GAT_882_gat), .Y(G2662GAT_882_ngat) );
INVXL U_g3089 (.A(G2659GAT_877_gat), .Y(G2659GAT_877_ngat) );
INVXL U_g3090 (.A(G2660GAT_884_gat), .Y(G2660GAT_884_ngat) );
INVXL U_g3091 (.A(G2657GAT_879_gat), .Y(G2657GAT_879_ngat) );
INVXL U_g3092 (.A(G2658GAT_885_gat), .Y(G2658GAT_885_ngat) );
INVXL U_g3093 (.A(G2655GAT_881_gat), .Y(G2655GAT_881_ngat) );
INVXL U_g3094 (.A(G2656GAT_886_gat), .Y(G2656GAT_886_ngat) );
INVXL U_g3095 (.A(G2653GAT_883_gat), .Y(G2653GAT_883_ngat) );
INVXL U_g3096 (.A(G2654GAT_887_gat), .Y(G2654GAT_887_ngat) );
INVXL U_g3097 (.A(G2743GAT_888_gat), .Y(G2743GAT_888_ngat) );
INVXL U_g3098 (.A(G2744GAT_889_gat), .Y(G2744GAT_889_ngat) );
INVXL U_g3099 (.A(G2739GAT_890_gat), .Y(G2739GAT_890_ngat) );
INVXL U_g3100 (.A(G2736GAT_891_gat), .Y(G2736GAT_891_ngat) );
INVXL U_g3101 (.A(G2733GAT_892_gat), .Y(G2733GAT_892_ngat) );
INVXL U_g3102 (.A(G2731GAT_893_gat), .Y(G2731GAT_893_ngat) );
INVXL U_g3103 (.A(G2732GAT_897_gat), .Y(G2732GAT_897_ngat) );
INVXL U_g3104 (.A(G2727GAT_899_gat), .Y(G2727GAT_899_ngat) );
INVXL U_g3105 (.A(G2724GAT_894_gat), .Y(G2724GAT_894_ngat) );
INVXL U_g3106 (.A(G1038GAT_122_gat), .Y(G1038GAT_122_ngat) );
INVXL U_g3107 (.A(G2721GAT_895_gat), .Y(G2721GAT_895_ngat) );
INVXL U_g3108 (.A(G990GAT_138_gat), .Y(G990GAT_138_ngat) );
INVXL U_g3109 (.A(G2718GAT_896_gat), .Y(G2718GAT_896_ngat) );
INVXL U_g3110 (.A(G942GAT_154_gat), .Y(G942GAT_154_ngat) );
INVXL U_g3111 (.A(G2715GAT_898_gat), .Y(G2715GAT_898_ngat) );
INVXL U_g3112 (.A(G894GAT_170_gat), .Y(G894GAT_170_ngat) );
INVXL U_g3113 (.A(G2712GAT_900_gat), .Y(G2712GAT_900_ngat) );
INVXL U_g3114 (.A(G846GAT_186_gat), .Y(G846GAT_186_ngat) );
INVXL U_g3115 (.A(G2709GAT_901_gat), .Y(G2709GAT_901_ngat) );
INVXL U_g3116 (.A(G798GAT_202_gat), .Y(G798GAT_202_ngat) );
INVXL U_g3117 (.A(G2706GAT_902_gat), .Y(G2706GAT_902_ngat) );
INVXL U_g3118 (.A(G750GAT_218_gat), .Y(G750GAT_218_ngat) );
INVXL U_g3119 (.A(G2703GAT_903_gat), .Y(G2703GAT_903_ngat) );
INVXL U_g3120 (.A(G702GAT_234_gat), .Y(G702GAT_234_ngat) );
INVXL U_g3121 (.A(G2700GAT_904_gat), .Y(G2700GAT_904_ngat) );
INVXL U_g3122 (.A(G654GAT_250_gat), .Y(G654GAT_250_ngat) );
INVXL U_g3123 (.A(G2697GAT_905_gat), .Y(G2697GAT_905_ngat) );
INVXL U_g3124 (.A(G606GAT_266_gat), .Y(G606GAT_266_ngat) );
INVXL U_g3125 (.A(G2694GAT_906_gat), .Y(G2694GAT_906_ngat) );
INVXL U_g3126 (.A(G558GAT_282_gat), .Y(G558GAT_282_ngat) );
INVXL U_g3127 (.A(G2801GAT_908_gat), .Y(G2801GAT_908_ngat) );
INVXL U_g3128 (.A(G2802GAT_909_gat), .Y(G2802GAT_909_ngat) );
INVXL U_g3129 (.A(G2797GAT_910_gat), .Y(G2797GAT_910_ngat) );
INVXL U_g3130 (.A(G2794GAT_911_gat), .Y(G2794GAT_911_ngat) );
INVXL U_g3131 (.A(G2791GAT_912_gat), .Y(G2791GAT_912_ngat) );
INVXL U_g3132 (.A(G2789GAT_913_gat), .Y(G2789GAT_913_ngat) );
INVXL U_g3133 (.A(G2790GAT_914_gat), .Y(G2790GAT_914_ngat) );
INVXL U_g3134 (.A(G2785GAT_915_gat), .Y(G2785GAT_915_ngat) );
INVXL U_g3135 (.A(G2803GAT_907_gat), .Y(G2803GAT_907_ngat) );
INVXL U_g3136 (.A(G1233GAT_57_gat), .Y(G1233GAT_57_ngat) );
INVXL U_g3137 (.A(G2781GAT_916_gat), .Y(G2781GAT_916_ngat) );
INVXL U_g3138 (.A(G2777GAT_917_gat), .Y(G2777GAT_917_ngat) );
INVXL U_g3139 (.A(G2773GAT_918_gat), .Y(G2773GAT_918_ngat) );
INVXL U_g3140 (.A(G2769GAT_919_gat), .Y(G2769GAT_919_ngat) );
INVXL U_g3141 (.A(G2765GAT_920_gat), .Y(G2765GAT_920_ngat) );
INVXL U_g3142 (.A(G2761GAT_921_gat), .Y(G2761GAT_921_ngat) );
INVXL U_g3143 (.A(G2757GAT_922_gat), .Y(G2757GAT_922_ngat) );
INVXL U_g3144 (.A(G2753GAT_923_gat), .Y(G2753GAT_923_ngat) );
INVXL U_g3145 (.A(G2749GAT_924_gat), .Y(G2749GAT_924_ngat) );
INVXL U_g3146 (.A(G2745GAT_925_gat), .Y(G2745GAT_925_ngat) );
INVXL U_g3147 (.A(G2873GAT_932_gat), .Y(G2873GAT_932_ngat) );
INVXL U_g3148 (.A(G2868GAT_927_gat), .Y(G2868GAT_927_ngat) );
INVXL U_g3149 (.A(G2869GAT_928_gat), .Y(G2869GAT_928_ngat) );
INVXL U_g3150 (.A(G2864GAT_929_gat), .Y(G2864GAT_929_ngat) );
INVXL U_g3151 (.A(G2861GAT_930_gat), .Y(G2861GAT_930_ngat) );
INVXL U_g3152 (.A(G2858GAT_936_gat), .Y(G2858GAT_936_ngat) );
INVXL U_g3153 (.A(G2856GAT_931_gat), .Y(G2856GAT_931_ngat) );
INVXL U_g3154 (.A(G2857GAT_938_gat), .Y(G2857GAT_938_ngat) );
INVXL U_g3155 (.A(G2851GAT_933_gat), .Y(G2851GAT_933_ngat) );
INVXL U_g3156 (.A(G2852GAT_941_gat), .Y(G2852GAT_941_ngat) );
INVXL U_g3157 (.A(G2870GAT_926_gat), .Y(G2870GAT_926_ngat) );
INVXL U_g3158 (.A(G1185GAT_73_gat), .Y(G1185GAT_73_ngat) );
INVXL U_g3159 (.A(G2846GAT_934_gat), .Y(G2846GAT_934_ngat) );
INVXL U_g3160 (.A(G2847GAT_944_gat), .Y(G2847GAT_944_ngat) );
INVXL U_g3161 (.A(G2841GAT_935_gat), .Y(G2841GAT_935_ngat) );
INVXL U_g3162 (.A(G2842GAT_947_gat), .Y(G2842GAT_947_ngat) );
INVXL U_g3163 (.A(G2836GAT_937_gat), .Y(G2836GAT_937_ngat) );
INVXL U_g3164 (.A(G2837GAT_950_gat), .Y(G2837GAT_950_ngat) );
INVXL U_g3165 (.A(G2831GAT_940_gat), .Y(G2831GAT_940_ngat) );
INVXL U_g3166 (.A(G2832GAT_953_gat), .Y(G2832GAT_953_ngat) );
INVXL U_g3167 (.A(G2826GAT_943_gat), .Y(G2826GAT_943_ngat) );
INVXL U_g3168 (.A(G2827GAT_956_gat), .Y(G2827GAT_956_ngat) );
INVXL U_g3169 (.A(G2821GAT_946_gat), .Y(G2821GAT_946_ngat) );
INVXL U_g3170 (.A(G2822GAT_958_gat), .Y(G2822GAT_958_ngat) );
INVXL U_g3171 (.A(G2816GAT_949_gat), .Y(G2816GAT_949_ngat) );
INVXL U_g3172 (.A(G2817GAT_960_gat), .Y(G2817GAT_960_ngat) );
INVXL U_g3173 (.A(G2811GAT_952_gat), .Y(G2811GAT_952_ngat) );
INVXL U_g3174 (.A(G2812GAT_962_gat), .Y(G2812GAT_962_ngat) );
INVXL U_g3175 (.A(G2806GAT_955_gat), .Y(G2806GAT_955_ngat) );
INVXL U_g3176 (.A(G2807GAT_964_gat), .Y(G2807GAT_964_ngat) );
INVXL U_g3177 (.A(G1281GAT_41_gat), .Y(G1281GAT_41_ngat) );
INVXL U_g3178 (.A(G2923GAT_965_gat), .Y(G2923GAT_965_ngat) );
INVXL U_g3179 (.A(G2921GAT_966_gat), .Y(G2921GAT_966_ngat) );
INVXL U_g3180 (.A(G2922GAT_972_gat), .Y(G2922GAT_972_ngat) );
INVXL U_g3181 (.A(G2917GAT_974_gat), .Y(G2917GAT_974_ngat) );
INVXL U_g3182 (.A(G2912GAT_968_gat), .Y(G2912GAT_968_ngat) );
INVXL U_g3183 (.A(G2913GAT_969_gat), .Y(G2913GAT_969_ngat) );
INVXL U_g3184 (.A(G2908GAT_970_gat), .Y(G2908GAT_970_ngat) );
INVXL U_g3185 (.A(G2914GAT_967_gat), .Y(G2914GAT_967_ngat) );
INVXL U_g3186 (.A(G1137GAT_89_gat), .Y(G1137GAT_89_ngat) );
INVXL U_g3187 (.A(G2905GAT_971_gat), .Y(G2905GAT_971_ngat) );
INVXL U_g3188 (.A(G2853GAT_939_gat), .Y(G2853GAT_939_ngat) );
INVXL U_g3189 (.A(G2902GAT_973_gat), .Y(G2902GAT_973_ngat) );
INVXL U_g3190 (.A(G2848GAT_942_gat), .Y(G2848GAT_942_ngat) );
INVXL U_g3191 (.A(G2899GAT_975_gat), .Y(G2899GAT_975_ngat) );
INVXL U_g3192 (.A(G2843GAT_945_gat), .Y(G2843GAT_945_ngat) );
INVXL U_g3193 (.A(G2896GAT_976_gat), .Y(G2896GAT_976_ngat) );
INVXL U_g3194 (.A(G2838GAT_948_gat), .Y(G2838GAT_948_ngat) );
INVXL U_g3195 (.A(G2893GAT_977_gat), .Y(G2893GAT_977_ngat) );
INVXL U_g3196 (.A(G2833GAT_951_gat), .Y(G2833GAT_951_ngat) );
INVXL U_g3197 (.A(G2890GAT_978_gat), .Y(G2890GAT_978_ngat) );
INVXL U_g3198 (.A(G2828GAT_954_gat), .Y(G2828GAT_954_ngat) );
INVXL U_g3199 (.A(G2887GAT_979_gat), .Y(G2887GAT_979_ngat) );
INVXL U_g3200 (.A(G2823GAT_957_gat), .Y(G2823GAT_957_ngat) );
INVXL U_g3201 (.A(G2884GAT_980_gat), .Y(G2884GAT_980_ngat) );
INVXL U_g3202 (.A(G2818GAT_959_gat), .Y(G2818GAT_959_ngat) );
INVXL U_g3203 (.A(G2881GAT_981_gat), .Y(G2881GAT_981_ngat) );
INVXL U_g3204 (.A(G2813GAT_961_gat), .Y(G2813GAT_961_ngat) );
INVXL U_g3205 (.A(G2878GAT_982_gat), .Y(G2878GAT_982_ngat) );
INVXL U_g3206 (.A(G2808GAT_963_gat), .Y(G2808GAT_963_ngat) );
INVXL U_g3207 (.A(G2983GAT_984_gat), .Y(G2983GAT_984_ngat) );
INVXL U_g3208 (.A(G2980GAT_985_gat), .Y(G2980GAT_985_ngat) );
INVXL U_g3209 (.A(G2977GAT_986_gat), .Y(G2977GAT_986_ngat) );
INVXL U_g3210 (.A(G2975GAT_987_gat), .Y(G2975GAT_987_ngat) );
INVXL U_g3211 (.A(G2976GAT_990_gat), .Y(G2976GAT_990_ngat) );
INVXL U_g3212 (.A(G2971GAT_991_gat), .Y(G2971GAT_991_ngat) );
INVXL U_g3213 (.A(G2966GAT_989_gat), .Y(G2966GAT_989_ngat) );
INVXL U_g3214 (.A(G2967GAT_992_gat), .Y(G2967GAT_992_ngat) );
INVXL U_g3215 (.A(G2962GAT_993_gat), .Y(G2962GAT_993_ngat) );
INVXL U_g3216 (.A(G2958GAT_994_gat), .Y(G2958GAT_994_ngat) );
INVXL U_g3217 (.A(G2954GAT_995_gat), .Y(G2954GAT_995_ngat) );
INVXL U_g3218 (.A(G2950GAT_996_gat), .Y(G2950GAT_996_ngat) );
INVXL U_g3219 (.A(G2968GAT_988_gat), .Y(G2968GAT_988_ngat) );
INVXL U_g3220 (.A(G1089GAT_105_gat), .Y(G1089GAT_105_ngat) );
INVXL U_g3221 (.A(G2946GAT_997_gat), .Y(G2946GAT_997_ngat) );
INVXL U_g3222 (.A(G2942GAT_998_gat), .Y(G2942GAT_998_ngat) );
INVXL U_g3223 (.A(G2938GAT_999_gat), .Y(G2938GAT_999_ngat) );
INVXL U_g3224 (.A(G2934GAT_1000_gat), .Y(G2934GAT_1000_ngat) );
INVXL U_g3225 (.A(G2930GAT_1001_gat), .Y(G2930GAT_1001_ngat) );
INVXL U_g3226 (.A(G2926GAT_1002_gat), .Y(G2926GAT_1002_ngat) );
INVXL U_g3227 (.A(G3026GAT_1003_gat), .Y(G3026GAT_1003_ngat) );
INVXL U_g3228 (.A(G3027GAT_1004_gat), .Y(G3027GAT_1004_ngat) );
INVXL U_g3229 (.A(G3022GAT_1005_gat), .Y(G3022GAT_1005_ngat) );
INVXL U_g3230 (.A(G3019GAT_1006_gat), .Y(G3019GAT_1006_ngat) );
INVXL U_g3231 (.A(G3016GAT_1007_gat), .Y(G3016GAT_1007_ngat) );
INVXL U_g3232 (.A(G3014GAT_1008_gat), .Y(G3014GAT_1008_ngat) );
INVXL U_g3233 (.A(G3015GAT_1013_gat), .Y(G3015GAT_1013_ngat) );
INVXL U_g3234 (.A(G3010GAT_1015_gat), .Y(G3010GAT_1015_ngat) );
INVXL U_g3235 (.A(G3005GAT_1010_gat), .Y(G3005GAT_1010_ngat) );
INVXL U_g3236 (.A(G3006GAT_1017_gat), .Y(G3006GAT_1017_ngat) );
INVXL U_g3237 (.A(G3003GAT_1011_gat), .Y(G3003GAT_1011_ngat) );
INVXL U_g3238 (.A(G3004GAT_1019_gat), .Y(G3004GAT_1019_ngat) );
INVXL U_g3239 (.A(G3001GAT_1012_gat), .Y(G3001GAT_1012_ngat) );
INVXL U_g3240 (.A(G3002GAT_1021_gat), .Y(G3002GAT_1021_ngat) );
INVXL U_g3241 (.A(G2999GAT_1014_gat), .Y(G2999GAT_1014_ngat) );
INVXL U_g3242 (.A(G3000GAT_1023_gat), .Y(G3000GAT_1023_ngat) );
INVXL U_g3243 (.A(G2997GAT_1016_gat), .Y(G2997GAT_1016_ngat) );
INVXL U_g3244 (.A(G2998GAT_1025_gat), .Y(G2998GAT_1025_ngat) );
INVXL U_g3245 (.A(G3007GAT_1009_gat), .Y(G3007GAT_1009_ngat) );
INVXL U_g3246 (.A(G1041GAT_121_gat), .Y(G1041GAT_121_ngat) );
INVXL U_g3247 (.A(G2995GAT_1018_gat), .Y(G2995GAT_1018_ngat) );
INVXL U_g3248 (.A(G2996GAT_1027_gat), .Y(G2996GAT_1027_ngat) );
INVXL U_g3249 (.A(G2993GAT_1020_gat), .Y(G2993GAT_1020_ngat) );
INVXL U_g3250 (.A(G2994GAT_1028_gat), .Y(G2994GAT_1028_ngat) );
INVXL U_g3251 (.A(G2991GAT_1022_gat), .Y(G2991GAT_1022_ngat) );
INVXL U_g3252 (.A(G2992GAT_1029_gat), .Y(G2992GAT_1029_ngat) );
INVXL U_g3253 (.A(G2989GAT_1024_gat), .Y(G2989GAT_1024_ngat) );
INVXL U_g3254 (.A(G2990GAT_1030_gat), .Y(G2990GAT_1030_ngat) );
INVXL U_g3255 (.A(G2987GAT_1026_gat), .Y(G2987GAT_1026_ngat) );
INVXL U_g3256 (.A(G2988GAT_1031_gat), .Y(G2988GAT_1031_ngat) );
INVXL U_g3257 (.A(G3074GAT_1033_gat), .Y(G3074GAT_1033_ngat) );
INVXL U_g3258 (.A(G3075GAT_1034_gat), .Y(G3075GAT_1034_ngat) );
INVXL U_g3259 (.A(G3070GAT_1035_gat), .Y(G3070GAT_1035_ngat) );
INVXL U_g3260 (.A(G3067GAT_1036_gat), .Y(G3067GAT_1036_ngat) );
INVXL U_g3261 (.A(G3064GAT_1037_gat), .Y(G3064GAT_1037_ngat) );
INVXL U_g3262 (.A(G3062GAT_1038_gat), .Y(G3062GAT_1038_ngat) );
INVXL U_g3263 (.A(G3063GAT_1043_gat), .Y(G3063GAT_1043_ngat) );
INVXL U_g3264 (.A(G3058GAT_1045_gat), .Y(G3058GAT_1045_ngat) );
INVXL U_g3265 (.A(G3076GAT_1032_gat), .Y(G3076GAT_1032_ngat) );
INVXL U_g3266 (.A(G1236GAT_56_gat), .Y(G1236GAT_56_ngat) );
INVXL U_g3267 (.A(G3055GAT_1039_gat), .Y(G3055GAT_1039_ngat) );
INVXL U_g3268 (.A(G993GAT_137_gat), .Y(G993GAT_137_ngat) );
INVXL U_g3269 (.A(G3052GAT_1040_gat), .Y(G3052GAT_1040_ngat) );
INVXL U_g3270 (.A(G945GAT_153_gat), .Y(G945GAT_153_ngat) );
INVXL U_g3271 (.A(G3049GAT_1041_gat), .Y(G3049GAT_1041_ngat) );
INVXL U_g3272 (.A(G897GAT_169_gat), .Y(G897GAT_169_ngat) );
INVXL U_g3273 (.A(G3046GAT_1042_gat), .Y(G3046GAT_1042_ngat) );
INVXL U_g3274 (.A(G849GAT_185_gat), .Y(G849GAT_185_ngat) );
INVXL U_g3275 (.A(G3043GAT_1044_gat), .Y(G3043GAT_1044_ngat) );
INVXL U_g3276 (.A(G801GAT_201_gat), .Y(G801GAT_201_ngat) );
INVXL U_g3277 (.A(G3040GAT_1046_gat), .Y(G3040GAT_1046_ngat) );
INVXL U_g3278 (.A(G753GAT_217_gat), .Y(G753GAT_217_ngat) );
INVXL U_g3279 (.A(G3037GAT_1047_gat), .Y(G3037GAT_1047_ngat) );
INVXL U_g3280 (.A(G705GAT_233_gat), .Y(G705GAT_233_ngat) );
INVXL U_g3281 (.A(G3034GAT_1048_gat), .Y(G3034GAT_1048_ngat) );
INVXL U_g3282 (.A(G657GAT_249_gat), .Y(G657GAT_249_ngat) );
INVXL U_g3283 (.A(G3031GAT_1049_gat), .Y(G3031GAT_1049_ngat) );
INVXL U_g3284 (.A(G609GAT_265_gat), .Y(G609GAT_265_ngat) );
INVXL U_g3285 (.A(G3028GAT_1050_gat), .Y(G3028GAT_1050_ngat) );
INVXL U_g3286 (.A(G561GAT_281_gat), .Y(G561GAT_281_ngat) );
INVXL U_g3287 (.A(G3136GAT_1058_gat), .Y(G3136GAT_1058_ngat) );
INVXL U_g3288 (.A(G3131GAT_1052_gat), .Y(G3131GAT_1052_ngat) );
INVXL U_g3289 (.A(G3132GAT_1053_gat), .Y(G3132GAT_1053_ngat) );
INVXL U_g3290 (.A(G3127GAT_1054_gat), .Y(G3127GAT_1054_ngat) );
INVXL U_g3291 (.A(G3124GAT_1055_gat), .Y(G3124GAT_1055_ngat) );
INVXL U_g3292 (.A(G3121GAT_1056_gat), .Y(G3121GAT_1056_ngat) );
INVXL U_g3293 (.A(G3119GAT_1057_gat), .Y(G3119GAT_1057_ngat) );
INVXL U_g3294 (.A(G3120GAT_1059_gat), .Y(G3120GAT_1059_ngat) );
INVXL U_g3295 (.A(G3115GAT_1060_gat), .Y(G3115GAT_1060_ngat) );
INVXL U_g3296 (.A(G3111GAT_1061_gat), .Y(G3111GAT_1061_ngat) );
INVXL U_g3297 (.A(G3133GAT_1051_gat), .Y(G3133GAT_1051_ngat) );
INVXL U_g3298 (.A(G1188GAT_72_gat), .Y(G1188GAT_72_ngat) );
INVXL U_g3299 (.A(G3107GAT_1062_gat), .Y(G3107GAT_1062_ngat) );
INVXL U_g3300 (.A(G3103GAT_1063_gat), .Y(G3103GAT_1063_ngat) );
INVXL U_g3301 (.A(G3099GAT_1064_gat), .Y(G3099GAT_1064_ngat) );
INVXL U_g3302 (.A(G3095GAT_1065_gat), .Y(G3095GAT_1065_ngat) );
INVXL U_g3303 (.A(G3091GAT_1066_gat), .Y(G3091GAT_1066_ngat) );
INVXL U_g3304 (.A(G3087GAT_1067_gat), .Y(G3087GAT_1067_ngat) );
INVXL U_g3305 (.A(G3083GAT_1068_gat), .Y(G3083GAT_1068_ngat) );
INVXL U_g3306 (.A(G3079GAT_1069_gat), .Y(G3079GAT_1069_ngat) );
INVXL U_g3307 (.A(G1284GAT_40_gat), .Y(G1284GAT_40_ngat) );
INVXL U_g3308 (.A(G3208GAT_1070_gat), .Y(G3208GAT_1070_ngat) );
INVXL U_g3309 (.A(G3206GAT_1071_gat), .Y(G3206GAT_1071_ngat) );
INVXL U_g3310 (.A(G3207GAT_1078_gat), .Y(G3207GAT_1078_ngat) );
INVXL U_g3311 (.A(G3202GAT_1080_gat), .Y(G3202GAT_1080_ngat) );
INVXL U_g3312 (.A(G3197GAT_1073_gat), .Y(G3197GAT_1073_ngat) );
INVXL U_g3313 (.A(G3198GAT_1074_gat), .Y(G3198GAT_1074_ngat) );
INVXL U_g3314 (.A(G3193GAT_1075_gat), .Y(G3193GAT_1075_ngat) );
INVXL U_g3315 (.A(G3190GAT_1076_gat), .Y(G3190GAT_1076_ngat) );
INVXL U_g3316 (.A(G3187GAT_1084_gat), .Y(G3187GAT_1084_ngat) );
INVXL U_g3317 (.A(G3185GAT_1077_gat), .Y(G3185GAT_1077_ngat) );
INVXL U_g3318 (.A(G3186GAT_1086_gat), .Y(G3186GAT_1086_ngat) );
INVXL U_g3319 (.A(G3180GAT_1079_gat), .Y(G3180GAT_1079_ngat) );
INVXL U_g3320 (.A(G3181GAT_1089_gat), .Y(G3181GAT_1089_ngat) );
INVXL U_g3321 (.A(G3175GAT_1081_gat), .Y(G3175GAT_1081_ngat) );
INVXL U_g3322 (.A(G3176GAT_1092_gat), .Y(G3176GAT_1092_ngat) );
INVXL U_g3323 (.A(G3199GAT_1072_gat), .Y(G3199GAT_1072_ngat) );
INVXL U_g3324 (.A(G1140GAT_88_gat), .Y(G1140GAT_88_ngat) );
INVXL U_g3325 (.A(G3170GAT_1082_gat), .Y(G3170GAT_1082_ngat) );
INVXL U_g3326 (.A(G3171GAT_1095_gat), .Y(G3171GAT_1095_ngat) );
INVXL U_g3327 (.A(G3165GAT_1083_gat), .Y(G3165GAT_1083_ngat) );
INVXL U_g3328 (.A(G3166GAT_1098_gat), .Y(G3166GAT_1098_ngat) );
INVXL U_g3329 (.A(G3160GAT_1085_gat), .Y(G3160GAT_1085_ngat) );
INVXL U_g3330 (.A(G3161GAT_1100_gat), .Y(G3161GAT_1100_ngat) );
INVXL U_g3331 (.A(G3155GAT_1088_gat), .Y(G3155GAT_1088_ngat) );
INVXL U_g3332 (.A(G3156GAT_1102_gat), .Y(G3156GAT_1102_ngat) );
INVXL U_g3333 (.A(G3150GAT_1091_gat), .Y(G3150GAT_1091_ngat) );
INVXL U_g3334 (.A(G3151GAT_1104_gat), .Y(G3151GAT_1104_ngat) );
INVXL U_g3335 (.A(G3145GAT_1094_gat), .Y(G3145GAT_1094_ngat) );
INVXL U_g3336 (.A(G3146GAT_1106_gat), .Y(G3146GAT_1106_ngat) );
INVXL U_g3337 (.A(G3140GAT_1097_gat), .Y(G3140GAT_1097_ngat) );
INVXL U_g3338 (.A(G3141GAT_1108_gat), .Y(G3141GAT_1108_ngat) );
INVXL U_g3339 (.A(G3260GAT_1109_gat), .Y(G3260GAT_1109_ngat) );
INVXL U_g3340 (.A(G3257GAT_1110_gat), .Y(G3257GAT_1110_ngat) );
INVXL U_g3341 (.A(G3254GAT_1111_gat), .Y(G3254GAT_1111_ngat) );
INVXL U_g3342 (.A(G3252GAT_1112_gat), .Y(G3252GAT_1112_ngat) );
INVXL U_g3343 (.A(G3253GAT_1119_gat), .Y(G3253GAT_1119_ngat) );
INVXL U_g3344 (.A(G3248GAT_1121_gat), .Y(G3248GAT_1121_ngat) );
INVXL U_g3345 (.A(G3243GAT_1114_gat), .Y(G3243GAT_1114_ngat) );
INVXL U_g3346 (.A(G3244GAT_1115_gat), .Y(G3244GAT_1115_ngat) );
INVXL U_g3347 (.A(G3239GAT_1116_gat), .Y(G3239GAT_1116_ngat) );
INVXL U_g3348 (.A(G3245GAT_1113_gat), .Y(G3245GAT_1113_ngat) );
INVXL U_g3349 (.A(G1092GAT_104_gat), .Y(G1092GAT_104_ngat) );
INVXL U_g3350 (.A(G3236GAT_1117_gat), .Y(G3236GAT_1117_ngat) );
INVXL U_g3351 (.A(G3182GAT_1087_gat), .Y(G3182GAT_1087_ngat) );
INVXL U_g3352 (.A(G3233GAT_1118_gat), .Y(G3233GAT_1118_ngat) );
INVXL U_g3353 (.A(G3177GAT_1090_gat), .Y(G3177GAT_1090_ngat) );
INVXL U_g3354 (.A(G3230GAT_1120_gat), .Y(G3230GAT_1120_ngat) );
INVXL U_g3355 (.A(G3172GAT_1093_gat), .Y(G3172GAT_1093_ngat) );
INVXL U_g3356 (.A(G3227GAT_1122_gat), .Y(G3227GAT_1122_ngat) );
INVXL U_g3357 (.A(G3167GAT_1096_gat), .Y(G3167GAT_1096_ngat) );
INVXL U_g3358 (.A(G3224GAT_1123_gat), .Y(G3224GAT_1123_ngat) );
INVXL U_g3359 (.A(G3162GAT_1099_gat), .Y(G3162GAT_1099_ngat) );
INVXL U_g3360 (.A(G3221GAT_1124_gat), .Y(G3221GAT_1124_ngat) );
INVXL U_g3361 (.A(G3157GAT_1101_gat), .Y(G3157GAT_1101_ngat) );
INVXL U_g3362 (.A(G3218GAT_1125_gat), .Y(G3218GAT_1125_ngat) );
INVXL U_g3363 (.A(G3152GAT_1103_gat), .Y(G3152GAT_1103_ngat) );
INVXL U_g3364 (.A(G3215GAT_1126_gat), .Y(G3215GAT_1126_ngat) );
INVXL U_g3365 (.A(G3147GAT_1105_gat), .Y(G3147GAT_1105_ngat) );
INVXL U_g3366 (.A(G3212GAT_1127_gat), .Y(G3212GAT_1127_ngat) );
INVXL U_g3367 (.A(G3142GAT_1107_gat), .Y(G3142GAT_1107_ngat) );
INVXL U_g3368 (.A(G3321GAT_1129_gat), .Y(G3321GAT_1129_ngat) );
INVXL U_g3369 (.A(G3322GAT_1130_gat), .Y(G3322GAT_1130_ngat) );
INVXL U_g3370 (.A(G3317GAT_1131_gat), .Y(G3317GAT_1131_ngat) );
INVXL U_g3371 (.A(G3314GAT_1132_gat), .Y(G3314GAT_1132_ngat) );
INVXL U_g3372 (.A(G3311GAT_1133_gat), .Y(G3311GAT_1133_ngat) );
INVXL U_g3373 (.A(G3309GAT_1134_gat), .Y(G3309GAT_1134_ngat) );
INVXL U_g3374 (.A(G3310GAT_1137_gat), .Y(G3310GAT_1137_ngat) );
INVXL U_g3375 (.A(G3305GAT_1138_gat), .Y(G3305GAT_1138_ngat) );
INVXL U_g3376 (.A(G3300GAT_1136_gat), .Y(G3300GAT_1136_ngat) );
INVXL U_g3377 (.A(G3301GAT_1139_gat), .Y(G3301GAT_1139_ngat) );
INVXL U_g3378 (.A(G3296GAT_1140_gat), .Y(G3296GAT_1140_ngat) );
INVXL U_g3379 (.A(G3292GAT_1141_gat), .Y(G3292GAT_1141_ngat) );
INVXL U_g3380 (.A(G3288GAT_1142_gat), .Y(G3288GAT_1142_ngat) );
INVXL U_g3381 (.A(G3284GAT_1143_gat), .Y(G3284GAT_1143_ngat) );
INVXL U_g3382 (.A(G3280GAT_1144_gat), .Y(G3280GAT_1144_ngat) );
INVXL U_g3383 (.A(G3302GAT_1135_gat), .Y(G3302GAT_1135_ngat) );
INVXL U_g3384 (.A(G1044GAT_120_gat), .Y(G1044GAT_120_ngat) );
INVXL U_g3385 (.A(G3276GAT_1145_gat), .Y(G3276GAT_1145_ngat) );
INVXL U_g3386 (.A(G3272GAT_1146_gat), .Y(G3272GAT_1146_ngat) );
INVXL U_g3387 (.A(G3268GAT_1147_gat), .Y(G3268GAT_1147_ngat) );
INVXL U_g3388 (.A(G3264GAT_1148_gat), .Y(G3264GAT_1148_ngat) );
INVXL U_g3389 (.A(G3360GAT_1150_gat), .Y(G3360GAT_1150_ngat) );
INVXL U_g3390 (.A(G3361GAT_1151_gat), .Y(G3361GAT_1151_ngat) );
INVXL U_g3391 (.A(G3356GAT_1152_gat), .Y(G3356GAT_1152_ngat) );
INVXL U_g3392 (.A(G3353GAT_1153_gat), .Y(G3353GAT_1153_ngat) );
INVXL U_g3393 (.A(G3350GAT_1154_gat), .Y(G3350GAT_1154_ngat) );
INVXL U_g3394 (.A(G3348GAT_1155_gat), .Y(G3348GAT_1155_ngat) );
INVXL U_g3395 (.A(G3349GAT_1161_gat), .Y(G3349GAT_1161_ngat) );
INVXL U_g3396 (.A(G3344GAT_1163_gat), .Y(G3344GAT_1163_ngat) );
INVXL U_g3397 (.A(G3339GAT_1157_gat), .Y(G3339GAT_1157_ngat) );
INVXL U_g3398 (.A(G3340GAT_1165_gat), .Y(G3340GAT_1165_ngat) );
INVXL U_g3399 (.A(G3362GAT_1149_gat), .Y(G3362GAT_1149_ngat) );
INVXL U_g3400 (.A(G1239GAT_55_gat), .Y(G1239GAT_55_ngat) );
INVXL U_g3401 (.A(G3337GAT_1158_gat), .Y(G3337GAT_1158_ngat) );
INVXL U_g3402 (.A(G3338GAT_1167_gat), .Y(G3338GAT_1167_ngat) );
INVXL U_g3403 (.A(G3335GAT_1159_gat), .Y(G3335GAT_1159_ngat) );
INVXL U_g3404 (.A(G3336GAT_1169_gat), .Y(G3336GAT_1169_ngat) );
INVXL U_g3405 (.A(G3333GAT_1160_gat), .Y(G3333GAT_1160_ngat) );
INVXL U_g3406 (.A(G3334GAT_1171_gat), .Y(G3334GAT_1171_ngat) );
INVXL U_g3407 (.A(G3331GAT_1162_gat), .Y(G3331GAT_1162_ngat) );
INVXL U_g3408 (.A(G3332GAT_1172_gat), .Y(G3332GAT_1172_ngat) );
INVXL U_g3409 (.A(G3329GAT_1164_gat), .Y(G3329GAT_1164_ngat) );
INVXL U_g3410 (.A(G3330GAT_1173_gat), .Y(G3330GAT_1173_ngat) );
INVXL U_g3411 (.A(G3341GAT_1156_gat), .Y(G3341GAT_1156_ngat) );
INVXL U_g3412 (.A(G996GAT_136_gat), .Y(G996GAT_136_ngat) );
INVXL U_g3413 (.A(G3327GAT_1166_gat), .Y(G3327GAT_1166_ngat) );
INVXL U_g3414 (.A(G3328GAT_1174_gat), .Y(G3328GAT_1174_ngat) );
INVXL U_g3415 (.A(G3325GAT_1168_gat), .Y(G3325GAT_1168_ngat) );
INVXL U_g3416 (.A(G3326GAT_1175_gat), .Y(G3326GAT_1175_ngat) );
INVXL U_g3417 (.A(G3323GAT_1170_gat), .Y(G3323GAT_1170_ngat) );
INVXL U_g3418 (.A(G3324GAT_1176_gat), .Y(G3324GAT_1176_ngat) );
INVXL U_g3419 (.A(G3413GAT_1185_gat), .Y(G3413GAT_1185_ngat) );
INVXL U_g3420 (.A(G3408GAT_1178_gat), .Y(G3408GAT_1178_ngat) );
INVXL U_g3421 (.A(G3409GAT_1179_gat), .Y(G3409GAT_1179_ngat) );
INVXL U_g3422 (.A(G3404GAT_1180_gat), .Y(G3404GAT_1180_ngat) );
INVXL U_g3423 (.A(G3401GAT_1181_gat), .Y(G3401GAT_1181_ngat) );
INVXL U_g3424 (.A(G3398GAT_1182_gat), .Y(G3398GAT_1182_ngat) );
INVXL U_g3425 (.A(G3396GAT_1183_gat), .Y(G3396GAT_1183_ngat) );
INVXL U_g3426 (.A(G3397GAT_1190_gat), .Y(G3397GAT_1190_ngat) );
INVXL U_g3427 (.A(G3392GAT_1192_gat), .Y(G3392GAT_1192_ngat) );
INVXL U_g3428 (.A(G3410GAT_1177_gat), .Y(G3410GAT_1177_ngat) );
INVXL U_g3429 (.A(G1191GAT_71_gat), .Y(G1191GAT_71_ngat) );
INVXL U_g3430 (.A(G3389GAT_1184_gat), .Y(G3389GAT_1184_ngat) );
INVXL U_g3431 (.A(G948GAT_152_gat), .Y(G948GAT_152_ngat) );
INVXL U_g3432 (.A(G3386GAT_1186_gat), .Y(G3386GAT_1186_ngat) );
INVXL U_g3433 (.A(G900GAT_168_gat), .Y(G900GAT_168_ngat) );
INVXL U_g3434 (.A(G3383GAT_1187_gat), .Y(G3383GAT_1187_ngat) );
INVXL U_g3435 (.A(G852GAT_184_gat), .Y(G852GAT_184_ngat) );
INVXL U_g3436 (.A(G3380GAT_1188_gat), .Y(G3380GAT_1188_ngat) );
INVXL U_g3437 (.A(G804GAT_200_gat), .Y(G804GAT_200_ngat) );
INVXL U_g3438 (.A(G3377GAT_1189_gat), .Y(G3377GAT_1189_ngat) );
INVXL U_g3439 (.A(G756GAT_216_gat), .Y(G756GAT_216_ngat) );
INVXL U_g3440 (.A(G3374GAT_1191_gat), .Y(G3374GAT_1191_ngat) );
INVXL U_g3441 (.A(G708GAT_232_gat), .Y(G708GAT_232_ngat) );
INVXL U_g3442 (.A(G3371GAT_1193_gat), .Y(G3371GAT_1193_ngat) );
INVXL U_g3443 (.A(G660GAT_248_gat), .Y(G660GAT_248_ngat) );
INVXL U_g3444 (.A(G3368GAT_1194_gat), .Y(G3368GAT_1194_ngat) );
INVXL U_g3445 (.A(G612GAT_264_gat), .Y(G612GAT_264_ngat) );
INVXL U_g3446 (.A(G3365GAT_1195_gat), .Y(G3365GAT_1195_ngat) );
INVXL U_g3447 (.A(G564GAT_280_gat), .Y(G564GAT_280_ngat) );
INVXL U_g3448 (.A(G1287GAT_39_gat), .Y(G1287GAT_39_ngat) );
INVXL U_g3449 (.A(G3476GAT_1196_gat), .Y(G3476GAT_1196_ngat) );
INVXL U_g3450 (.A(G3474GAT_1197_gat), .Y(G3474GAT_1197_ngat) );
INVXL U_g3451 (.A(G3475GAT_1205_gat), .Y(G3475GAT_1205_ngat) );
INVXL U_g3452 (.A(G3470GAT_1206_gat), .Y(G3470GAT_1206_ngat) );
INVXL U_g3453 (.A(G3465GAT_1199_gat), .Y(G3465GAT_1199_ngat) );
INVXL U_g3454 (.A(G3466GAT_1200_gat), .Y(G3466GAT_1200_ngat) );
INVXL U_g3455 (.A(G3461GAT_1201_gat), .Y(G3461GAT_1201_ngat) );
INVXL U_g3456 (.A(G3458GAT_1202_gat), .Y(G3458GAT_1202_ngat) );
INVXL U_g3457 (.A(G3455GAT_1203_gat), .Y(G3455GAT_1203_ngat) );
INVXL U_g3458 (.A(G3453GAT_1204_gat), .Y(G3453GAT_1204_ngat) );
INVXL U_g3459 (.A(G3454GAT_1207_gat), .Y(G3454GAT_1207_ngat) );
INVXL U_g3460 (.A(G3449GAT_1208_gat), .Y(G3449GAT_1208_ngat) );
INVXL U_g3461 (.A(G3445GAT_1209_gat), .Y(G3445GAT_1209_ngat) );
INVXL U_g3462 (.A(G3441GAT_1210_gat), .Y(G3441GAT_1210_ngat) );
INVXL U_g3463 (.A(G3467GAT_1198_gat), .Y(G3467GAT_1198_ngat) );
INVXL U_g3464 (.A(G1143GAT_87_gat), .Y(G1143GAT_87_ngat) );
INVXL U_g3465 (.A(G3437GAT_1211_gat), .Y(G3437GAT_1211_ngat) );
INVXL U_g3466 (.A(G3433GAT_1212_gat), .Y(G3433GAT_1212_ngat) );
INVXL U_g3467 (.A(G3429GAT_1213_gat), .Y(G3429GAT_1213_ngat) );
INVXL U_g3468 (.A(G3425GAT_1214_gat), .Y(G3425GAT_1214_ngat) );
INVXL U_g3469 (.A(G3421GAT_1215_gat), .Y(G3421GAT_1215_ngat) );
INVXL U_g3470 (.A(G3417GAT_1216_gat), .Y(G3417GAT_1216_ngat) );
INVXL U_g3471 (.A(G3548GAT_1217_gat), .Y(G3548GAT_1217_ngat) );
INVXL U_g3472 (.A(G3545GAT_1218_gat), .Y(G3545GAT_1218_ngat) );
INVXL U_g3473 (.A(G3542GAT_1219_gat), .Y(G3542GAT_1219_ngat) );
INVXL U_g3474 (.A(G3540GAT_1220_gat), .Y(G3540GAT_1220_ngat) );
INVXL U_g3475 (.A(G3541GAT_1228_gat), .Y(G3541GAT_1228_ngat) );
INVXL U_g3476 (.A(G3536GAT_1230_gat), .Y(G3536GAT_1230_ngat) );
INVXL U_g3477 (.A(G3531GAT_1222_gat), .Y(G3531GAT_1222_ngat) );
INVXL U_g3478 (.A(G3532GAT_1223_gat), .Y(G3532GAT_1223_ngat) );
INVXL U_g3479 (.A(G3527GAT_1224_gat), .Y(G3527GAT_1224_ngat) );
INVXL U_g3480 (.A(G3524GAT_1225_gat), .Y(G3524GAT_1225_ngat) );
INVXL U_g3481 (.A(G3521GAT_1234_gat), .Y(G3521GAT_1234_ngat) );
INVXL U_g3482 (.A(G3519GAT_1226_gat), .Y(G3519GAT_1226_ngat) );
INVXL U_g3483 (.A(G3520GAT_1236_gat), .Y(G3520GAT_1236_ngat) );
INVXL U_g3484 (.A(G3514GAT_1227_gat), .Y(G3514GAT_1227_ngat) );
INVXL U_g3485 (.A(G3515GAT_1239_gat), .Y(G3515GAT_1239_ngat) );
INVXL U_g3486 (.A(G3509GAT_1229_gat), .Y(G3509GAT_1229_ngat) );
INVXL U_g3487 (.A(G3510GAT_1242_gat), .Y(G3510GAT_1242_ngat) );
INVXL U_g3488 (.A(G3504GAT_1231_gat), .Y(G3504GAT_1231_ngat) );
INVXL U_g3489 (.A(G3505GAT_1244_gat), .Y(G3505GAT_1244_ngat) );
INVXL U_g3490 (.A(G3533GAT_1221_gat), .Y(G3533GAT_1221_ngat) );
INVXL U_g3491 (.A(G1095GAT_103_gat), .Y(G1095GAT_103_ngat) );
INVXL U_g3492 (.A(G3499GAT_1232_gat), .Y(G3499GAT_1232_ngat) );
INVXL U_g3493 (.A(G3500GAT_1246_gat), .Y(G3500GAT_1246_ngat) );
INVXL U_g3494 (.A(G3494GAT_1233_gat), .Y(G3494GAT_1233_ngat) );
INVXL U_g3495 (.A(G3495GAT_1248_gat), .Y(G3495GAT_1248_ngat) );
INVXL U_g3496 (.A(G3489GAT_1235_gat), .Y(G3489GAT_1235_ngat) );
INVXL U_g3497 (.A(G3490GAT_1250_gat), .Y(G3490GAT_1250_ngat) );
INVXL U_g3498 (.A(G3484GAT_1238_gat), .Y(G3484GAT_1238_ngat) );
INVXL U_g3499 (.A(G3485GAT_1252_gat), .Y(G3485GAT_1252_ngat) );
INVXL U_g3500 (.A(G3479GAT_1241_gat), .Y(G3479GAT_1241_ngat) );
INVXL U_g3501 (.A(G3480GAT_1254_gat), .Y(G3480GAT_1254_ngat) );
INVXL U_g3502 (.A(G3602GAT_1255_gat), .Y(G3602GAT_1255_ngat) );
INVXL U_g3503 (.A(G3603GAT_1256_gat), .Y(G3603GAT_1256_ngat) );
INVXL U_g3504 (.A(G3598GAT_1257_gat), .Y(G3598GAT_1257_ngat) );
INVXL U_g3505 (.A(G3595GAT_1258_gat), .Y(G3595GAT_1258_ngat) );
INVXL U_g3506 (.A(G3592GAT_1259_gat), .Y(G3592GAT_1259_ngat) );
INVXL U_g3507 (.A(G3590GAT_1260_gat), .Y(G3590GAT_1260_ngat) );
INVXL U_g3508 (.A(G3591GAT_1268_gat), .Y(G3591GAT_1268_ngat) );
INVXL U_g3509 (.A(G3586GAT_1270_gat), .Y(G3586GAT_1270_ngat) );
INVXL U_g3510 (.A(G3581GAT_1262_gat), .Y(G3581GAT_1262_ngat) );
INVXL U_g3511 (.A(G3582GAT_1263_gat), .Y(G3582GAT_1263_ngat) );
INVXL U_g3512 (.A(G3577GAT_1264_gat), .Y(G3577GAT_1264_ngat) );
INVXL U_g3513 (.A(G3583GAT_1261_gat), .Y(G3583GAT_1261_ngat) );
INVXL U_g3514 (.A(G1047GAT_119_gat), .Y(G1047GAT_119_ngat) );
INVXL U_g3515 (.A(G3574GAT_1265_gat), .Y(G3574GAT_1265_ngat) );
INVXL U_g3516 (.A(G3516GAT_1237_gat), .Y(G3516GAT_1237_ngat) );
INVXL U_g3517 (.A(G3571GAT_1266_gat), .Y(G3571GAT_1266_ngat) );
INVXL U_g3518 (.A(G3511GAT_1240_gat), .Y(G3511GAT_1240_ngat) );
INVXL U_g3519 (.A(G3568GAT_1267_gat), .Y(G3568GAT_1267_ngat) );
INVXL U_g3520 (.A(G3506GAT_1243_gat), .Y(G3506GAT_1243_ngat) );
INVXL U_g3521 (.A(G3565GAT_1269_gat), .Y(G3565GAT_1269_ngat) );
INVXL U_g3522 (.A(G3501GAT_1245_gat), .Y(G3501GAT_1245_ngat) );
INVXL U_g3523 (.A(G3562GAT_1271_gat), .Y(G3562GAT_1271_ngat) );
INVXL U_g3524 (.A(G3496GAT_1247_gat), .Y(G3496GAT_1247_ngat) );
INVXL U_g3525 (.A(G3559GAT_1272_gat), .Y(G3559GAT_1272_ngat) );
INVXL U_g3526 (.A(G3491GAT_1249_gat), .Y(G3491GAT_1249_ngat) );
INVXL U_g3527 (.A(G3556GAT_1273_gat), .Y(G3556GAT_1273_ngat) );
INVXL U_g3528 (.A(G3486GAT_1251_gat), .Y(G3486GAT_1251_ngat) );
INVXL U_g3529 (.A(G3553GAT_1274_gat), .Y(G3553GAT_1274_ngat) );
INVXL U_g3530 (.A(G3481GAT_1253_gat), .Y(G3481GAT_1253_ngat) );
INVXL U_g3531 (.A(G3657GAT_1277_gat), .Y(G3657GAT_1277_ngat) );
INVXL U_g3532 (.A(G3658GAT_1278_gat), .Y(G3658GAT_1278_ngat) );
INVXL U_g3533 (.A(G3653GAT_1279_gat), .Y(G3653GAT_1279_ngat) );
INVXL U_g3534 (.A(G3650GAT_1280_gat), .Y(G3650GAT_1280_ngat) );
INVXL U_g3535 (.A(G3647GAT_1281_gat), .Y(G3647GAT_1281_ngat) );
INVXL U_g3536 (.A(G3645GAT_1282_gat), .Y(G3645GAT_1282_ngat) );
INVXL U_g3537 (.A(G3646GAT_1285_gat), .Y(G3646GAT_1285_ngat) );
INVXL U_g3538 (.A(G3641GAT_1286_gat), .Y(G3641GAT_1286_ngat) );
INVXL U_g3539 (.A(G3636GAT_1284_gat), .Y(G3636GAT_1284_ngat) );
INVXL U_g3540 (.A(G3637GAT_1287_gat), .Y(G3637GAT_1287_ngat) );
INVXL U_g3541 (.A(G3632GAT_1288_gat), .Y(G3632GAT_1288_ngat) );
INVXL U_g3542 (.A(G3659GAT_1276_gat), .Y(G3659GAT_1276_ngat) );
INVXL U_g3543 (.A(G1242GAT_54_gat), .Y(G1242GAT_54_ngat) );
INVXL U_g3544 (.A(G3628GAT_1289_gat), .Y(G3628GAT_1289_ngat) );
INVXL U_g3545 (.A(G3624GAT_1290_gat), .Y(G3624GAT_1290_ngat) );
INVXL U_g3546 (.A(G3620GAT_1291_gat), .Y(G3620GAT_1291_ngat) );
INVXL U_g3547 (.A(G3616GAT_1292_gat), .Y(G3616GAT_1292_ngat) );
INVXL U_g3548 (.A(G3612GAT_1293_gat), .Y(G3612GAT_1293_ngat) );
INVXL U_g3549 (.A(G3638GAT_1283_gat), .Y(G3638GAT_1283_ngat) );
INVXL U_g3550 (.A(G999GAT_135_gat), .Y(G999GAT_135_ngat) );
INVXL U_g3551 (.A(G3608GAT_1294_gat), .Y(G3608GAT_1294_ngat) );
INVXL U_g3552 (.A(G3604GAT_1295_gat), .Y(G3604GAT_1295_ngat) );
INVXL U_g3553 (.A(G3702GAT_1305_gat), .Y(G3702GAT_1305_ngat) );
INVXL U_g3554 (.A(G3697GAT_1297_gat), .Y(G3697GAT_1297_ngat) );
INVXL U_g3555 (.A(G3698GAT_1298_gat), .Y(G3698GAT_1298_ngat) );
INVXL U_g3556 (.A(G3693GAT_1299_gat), .Y(G3693GAT_1299_ngat) );
INVXL U_g3557 (.A(G3690GAT_1300_gat), .Y(G3690GAT_1300_ngat) );
INVXL U_g3558 (.A(G3687GAT_1301_gat), .Y(G3687GAT_1301_ngat) );
INVXL U_g3559 (.A(G3685GAT_1302_gat), .Y(G3685GAT_1302_ngat) );
INVXL U_g3560 (.A(G3686GAT_1310_gat), .Y(G3686GAT_1310_ngat) );
INVXL U_g3561 (.A(G3681GAT_1312_gat), .Y(G3681GAT_1312_ngat) );
INVXL U_g3562 (.A(G3676GAT_1304_gat), .Y(G3676GAT_1304_ngat) );
INVXL U_g3563 (.A(G3677GAT_1314_gat), .Y(G3677GAT_1314_ngat) );
INVXL U_g3564 (.A(G3674GAT_1306_gat), .Y(G3674GAT_1306_ngat) );
INVXL U_g3565 (.A(G3675GAT_1316_gat), .Y(G3675GAT_1316_ngat) );
INVXL U_g3566 (.A(G3699GAT_1296_gat), .Y(G3699GAT_1296_ngat) );
INVXL U_g3567 (.A(G1194GAT_70_gat), .Y(G1194GAT_70_ngat) );
INVXL U_g3568 (.A(G3672GAT_1307_gat), .Y(G3672GAT_1307_ngat) );
INVXL U_g3569 (.A(G3673GAT_1317_gat), .Y(G3673GAT_1317_ngat) );
INVXL U_g3570 (.A(G3670GAT_1308_gat), .Y(G3670GAT_1308_ngat) );
INVXL U_g3571 (.A(G3671GAT_1318_gat), .Y(G3671GAT_1318_ngat) );
INVXL U_g3572 (.A(G3668GAT_1309_gat), .Y(G3668GAT_1309_ngat) );
INVXL U_g3573 (.A(G3669GAT_1319_gat), .Y(G3669GAT_1319_ngat) );
INVXL U_g3574 (.A(G3666GAT_1311_gat), .Y(G3666GAT_1311_ngat) );
INVXL U_g3575 (.A(G3667GAT_1320_gat), .Y(G3667GAT_1320_ngat) );
INVXL U_g3576 (.A(G3664GAT_1313_gat), .Y(G3664GAT_1313_ngat) );
INVXL U_g3577 (.A(G3665GAT_1321_gat), .Y(G3665GAT_1321_ngat) );
INVXL U_g3578 (.A(G3678GAT_1303_gat), .Y(G3678GAT_1303_ngat) );
INVXL U_g3579 (.A(G951GAT_151_gat), .Y(G951GAT_151_ngat) );
INVXL U_g3580 (.A(G3662GAT_1315_gat), .Y(G3662GAT_1315_ngat) );
INVXL U_g3581 (.A(G3663GAT_1322_gat), .Y(G3663GAT_1322_ngat) );
INVXL U_g3582 (.A(G1290GAT_38_gat), .Y(G1290GAT_38_ngat) );
INVXL U_g3583 (.A(G3757GAT_1323_gat), .Y(G3757GAT_1323_ngat) );
INVXL U_g3584 (.A(G3755GAT_1324_gat), .Y(G3755GAT_1324_ngat) );
INVXL U_g3585 (.A(G3756GAT_1333_gat), .Y(G3756GAT_1333_ngat) );
INVXL U_g3586 (.A(G3751GAT_1335_gat), .Y(G3751GAT_1335_ngat) );
INVXL U_g3587 (.A(G3746GAT_1326_gat), .Y(G3746GAT_1326_ngat) );
INVXL U_g3588 (.A(G3747GAT_1327_gat), .Y(G3747GAT_1327_ngat) );
INVXL U_g3589 (.A(G3742GAT_1328_gat), .Y(G3742GAT_1328_ngat) );
INVXL U_g3590 (.A(G3739GAT_1329_gat), .Y(G3739GAT_1329_ngat) );
INVXL U_g3591 (.A(G3736GAT_1330_gat), .Y(G3736GAT_1330_ngat) );
INVXL U_g3592 (.A(G3734GAT_1331_gat), .Y(G3734GAT_1331_ngat) );
INVXL U_g3593 (.A(G3735GAT_1340_gat), .Y(G3735GAT_1340_ngat) );
INVXL U_g3594 (.A(G3730GAT_1342_gat), .Y(G3730GAT_1342_ngat) );
INVXL U_g3595 (.A(G3748GAT_1325_gat), .Y(G3748GAT_1325_ngat) );
INVXL U_g3596 (.A(G1146GAT_86_gat), .Y(G1146GAT_86_ngat) );
INVXL U_g3597 (.A(G3727GAT_1332_gat), .Y(G3727GAT_1332_ngat) );
INVXL U_g3598 (.A(G903GAT_167_gat), .Y(G903GAT_167_ngat) );
INVXL U_g3599 (.A(G3724GAT_1334_gat), .Y(G3724GAT_1334_ngat) );
INVXL U_g3600 (.A(G855GAT_183_gat), .Y(G855GAT_183_ngat) );
INVXL U_g3601 (.A(G3721GAT_1336_gat), .Y(G3721GAT_1336_ngat) );
INVXL U_g3602 (.A(G807GAT_199_gat), .Y(G807GAT_199_ngat) );
INVXL U_g3603 (.A(G3718GAT_1337_gat), .Y(G3718GAT_1337_ngat) );
INVXL U_g3604 (.A(G759GAT_215_gat), .Y(G759GAT_215_ngat) );
INVXL U_g3605 (.A(G3715GAT_1338_gat), .Y(G3715GAT_1338_ngat) );
INVXL U_g3606 (.A(G711GAT_231_gat), .Y(G711GAT_231_ngat) );
INVXL U_g3607 (.A(G3712GAT_1339_gat), .Y(G3712GAT_1339_ngat) );
INVXL U_g3608 (.A(G663GAT_247_gat), .Y(G663GAT_247_ngat) );
INVXL U_g3609 (.A(G3709GAT_1341_gat), .Y(G3709GAT_1341_ngat) );
INVXL U_g3610 (.A(G615GAT_263_gat), .Y(G615GAT_263_ngat) );
INVXL U_g3611 (.A(G3706GAT_1343_gat), .Y(G3706GAT_1343_ngat) );
INVXL U_g3612 (.A(G567GAT_279_gat), .Y(G567GAT_279_ngat) );
INVXL U_g3613 (.A(G3821GAT_1344_gat), .Y(G3821GAT_1344_ngat) );
INVXL U_g3614 (.A(G3818GAT_1345_gat), .Y(G3818GAT_1345_ngat) );
INVXL U_g3615 (.A(G3815GAT_1346_gat), .Y(G3815GAT_1346_ngat) );
INVXL U_g3616 (.A(G3813GAT_1347_gat), .Y(G3813GAT_1347_ngat) );
INVXL U_g3617 (.A(G3814GAT_1355_gat), .Y(G3814GAT_1355_ngat) );
INVXL U_g3618 (.A(G3809GAT_1356_gat), .Y(G3809GAT_1356_ngat) );
INVXL U_g3619 (.A(G3804GAT_1349_gat), .Y(G3804GAT_1349_ngat) );
INVXL U_g3620 (.A(G3805GAT_1350_gat), .Y(G3805GAT_1350_ngat) );
INVXL U_g3621 (.A(G3800GAT_1351_gat), .Y(G3800GAT_1351_ngat) );
INVXL U_g3622 (.A(G3797GAT_1352_gat), .Y(G3797GAT_1352_ngat) );
INVXL U_g3623 (.A(G3794GAT_1353_gat), .Y(G3794GAT_1353_ngat) );
INVXL U_g3624 (.A(G3792GAT_1354_gat), .Y(G3792GAT_1354_ngat) );
INVXL U_g3625 (.A(G3793GAT_1357_gat), .Y(G3793GAT_1357_ngat) );
INVXL U_g3626 (.A(G3788GAT_1358_gat), .Y(G3788GAT_1358_ngat) );
INVXL U_g3627 (.A(G3784GAT_1359_gat), .Y(G3784GAT_1359_ngat) );
INVXL U_g3628 (.A(G3780GAT_1360_gat), .Y(G3780GAT_1360_ngat) );
INVXL U_g3629 (.A(G3776GAT_1361_gat), .Y(G3776GAT_1361_ngat) );
INVXL U_g3630 (.A(G3806GAT_1348_gat), .Y(G3806GAT_1348_ngat) );
INVXL U_g3631 (.A(G1098GAT_102_gat), .Y(G1098GAT_102_ngat) );
INVXL U_g3632 (.A(G3772GAT_1362_gat), .Y(G3772GAT_1362_ngat) );
INVXL U_g3633 (.A(G3768GAT_1363_gat), .Y(G3768GAT_1363_ngat) );
INVXL U_g3634 (.A(G3764GAT_1364_gat), .Y(G3764GAT_1364_ngat) );
INVXL U_g3635 (.A(G3760GAT_1365_gat), .Y(G3760GAT_1365_ngat) );
INVXL U_g3636 (.A(G3893GAT_1366_gat), .Y(G3893GAT_1366_ngat) );
INVXL U_g3637 (.A(G3894GAT_1367_gat), .Y(G3894GAT_1367_ngat) );
INVXL U_g3638 (.A(G3889GAT_1368_gat), .Y(G3889GAT_1368_ngat) );
INVXL U_g3639 (.A(G3886GAT_1369_gat), .Y(G3886GAT_1369_ngat) );
INVXL U_g3640 (.A(G3883GAT_1370_gat), .Y(G3883GAT_1370_ngat) );
INVXL U_g3641 (.A(G3881GAT_1371_gat), .Y(G3881GAT_1371_ngat) );
INVXL U_g3642 (.A(G3882GAT_1380_gat), .Y(G3882GAT_1380_ngat) );
INVXL U_g3643 (.A(G3877GAT_1382_gat), .Y(G3877GAT_1382_ngat) );
INVXL U_g3644 (.A(G3872GAT_1373_gat), .Y(G3872GAT_1373_ngat) );
INVXL U_g3645 (.A(G3873GAT_1374_gat), .Y(G3873GAT_1374_ngat) );
INVXL U_g3646 (.A(G3868GAT_1375_gat), .Y(G3868GAT_1375_ngat) );
INVXL U_g3647 (.A(G3865GAT_1376_gat), .Y(G3865GAT_1376_ngat) );
INVXL U_g3648 (.A(G3862GAT_1386_gat), .Y(G3862GAT_1386_ngat) );
INVXL U_g3649 (.A(G3860GAT_1377_gat), .Y(G3860GAT_1377_ngat) );
INVXL U_g3650 (.A(G3861GAT_1388_gat), .Y(G3861GAT_1388_ngat) );
INVXL U_g3651 (.A(G3855GAT_1378_gat), .Y(G3855GAT_1378_ngat) );
INVXL U_g3652 (.A(G3856GAT_1390_gat), .Y(G3856GAT_1390_ngat) );
INVXL U_g3653 (.A(G3850GAT_1379_gat), .Y(G3850GAT_1379_ngat) );
INVXL U_g3654 (.A(G3851GAT_1392_gat), .Y(G3851GAT_1392_ngat) );
INVXL U_g3655 (.A(G3845GAT_1381_gat), .Y(G3845GAT_1381_ngat) );
INVXL U_g3656 (.A(G3846GAT_1394_gat), .Y(G3846GAT_1394_ngat) );
INVXL U_g3657 (.A(G3840GAT_1383_gat), .Y(G3840GAT_1383_ngat) );
INVXL U_g3658 (.A(G3841GAT_1396_gat), .Y(G3841GAT_1396_ngat) );
INVXL U_g3659 (.A(G3874GAT_1372_gat), .Y(G3874GAT_1372_ngat) );
INVXL U_g3660 (.A(G1050GAT_118_gat), .Y(G1050GAT_118_ngat) );
INVXL U_g3661 (.A(G3835GAT_1384_gat), .Y(G3835GAT_1384_ngat) );
INVXL U_g3662 (.A(G3836GAT_1398_gat), .Y(G3836GAT_1398_ngat) );
INVXL U_g3663 (.A(G3830GAT_1385_gat), .Y(G3830GAT_1385_ngat) );
INVXL U_g3664 (.A(G3831GAT_1400_gat), .Y(G3831GAT_1400_ngat) );
INVXL U_g3665 (.A(G3825GAT_1387_gat), .Y(G3825GAT_1387_ngat) );
INVXL U_g3666 (.A(G3826GAT_1402_gat), .Y(G3826GAT_1402_ngat) );
INVXL U_g3667 (.A(G3942GAT_1404_gat), .Y(G3942GAT_1404_ngat) );
INVXL U_g3668 (.A(G3943GAT_1405_gat), .Y(G3943GAT_1405_ngat) );
INVXL U_g3669 (.A(G3938GAT_1406_gat), .Y(G3938GAT_1406_ngat) );
INVXL U_g3670 (.A(G3935GAT_1407_gat), .Y(G3935GAT_1407_ngat) );
INVXL U_g3671 (.A(G3932GAT_1408_gat), .Y(G3932GAT_1408_ngat) );
INVXL U_g3672 (.A(G3930GAT_1409_gat), .Y(G3930GAT_1409_ngat) );
INVXL U_g3673 (.A(G3931GAT_1418_gat), .Y(G3931GAT_1418_ngat) );
INVXL U_g3674 (.A(G3926GAT_1420_gat), .Y(G3926GAT_1420_ngat) );
INVXL U_g3675 (.A(G3921GAT_1411_gat), .Y(G3921GAT_1411_ngat) );
INVXL U_g3676 (.A(G3922GAT_1412_gat), .Y(G3922GAT_1412_ngat) );
INVXL U_g3677 (.A(G3917GAT_1413_gat), .Y(G3917GAT_1413_ngat) );
INVXL U_g3678 (.A(G3944GAT_1403_gat), .Y(G3944GAT_1403_ngat) );
INVXL U_g3679 (.A(G1245GAT_53_gat), .Y(G1245GAT_53_ngat) );
INVXL U_g3680 (.A(G3923GAT_1410_gat), .Y(G3923GAT_1410_ngat) );
INVXL U_g3681 (.A(G1002GAT_134_gat), .Y(G1002GAT_134_ngat) );
INVXL U_g3682 (.A(G3914GAT_1414_gat), .Y(G3914GAT_1414_ngat) );
INVXL U_g3683 (.A(G3857GAT_1389_gat), .Y(G3857GAT_1389_ngat) );
INVXL U_g3684 (.A(G3911GAT_1415_gat), .Y(G3911GAT_1415_ngat) );
INVXL U_g3685 (.A(G3852GAT_1391_gat), .Y(G3852GAT_1391_ngat) );
INVXL U_g3686 (.A(G3908GAT_1416_gat), .Y(G3908GAT_1416_ngat) );
INVXL U_g3687 (.A(G3847GAT_1393_gat), .Y(G3847GAT_1393_ngat) );
INVXL U_g3688 (.A(G3905GAT_1417_gat), .Y(G3905GAT_1417_ngat) );
INVXL U_g3689 (.A(G3842GAT_1395_gat), .Y(G3842GAT_1395_ngat) );
INVXL U_g3690 (.A(G3902GAT_1419_gat), .Y(G3902GAT_1419_ngat) );
INVXL U_g3691 (.A(G3837GAT_1397_gat), .Y(G3837GAT_1397_ngat) );
INVXL U_g3692 (.A(G3899GAT_1421_gat), .Y(G3899GAT_1421_ngat) );
INVXL U_g3693 (.A(G3832GAT_1399_gat), .Y(G3832GAT_1399_ngat) );
INVXL U_g3694 (.A(G3896GAT_1422_gat), .Y(G3896GAT_1422_ngat) );
INVXL U_g3695 (.A(G3827GAT_1401_gat), .Y(G3827GAT_1401_ngat) );
INVXL U_g3696 (.A(G4001GAT_1433_gat), .Y(G4001GAT_1433_ngat) );
INVXL U_g3697 (.A(G3996GAT_1425_gat), .Y(G3996GAT_1425_ngat) );
INVXL U_g3698 (.A(G3997GAT_1426_gat), .Y(G3997GAT_1426_ngat) );
INVXL U_g3699 (.A(G3992GAT_1427_gat), .Y(G3992GAT_1427_ngat) );
INVXL U_g3700 (.A(G3989GAT_1428_gat), .Y(G3989GAT_1428_ngat) );
INVXL U_g3701 (.A(G3986GAT_1429_gat), .Y(G3986GAT_1429_ngat) );
INVXL U_g3702 (.A(G3984GAT_1430_gat), .Y(G3984GAT_1430_ngat) );
INVXL U_g3703 (.A(G3985GAT_1434_gat), .Y(G3985GAT_1434_ngat) );
INVXL U_g3704 (.A(G3980GAT_1435_gat), .Y(G3980GAT_1435_ngat) );
INVXL U_g3705 (.A(G3975GAT_1432_gat), .Y(G3975GAT_1432_ngat) );
INVXL U_g3706 (.A(G3976GAT_1436_gat), .Y(G3976GAT_1436_ngat) );
INVXL U_g3707 (.A(G3971GAT_1437_gat), .Y(G3971GAT_1437_ngat) );
INVXL U_g3708 (.A(G3967GAT_1438_gat), .Y(G3967GAT_1438_ngat) );
INVXL U_g3709 (.A(G3998GAT_1424_gat), .Y(G3998GAT_1424_ngat) );
INVXL U_g3710 (.A(G1197GAT_69_gat), .Y(G1197GAT_69_ngat) );
INVXL U_g3711 (.A(G3963GAT_1439_gat), .Y(G3963GAT_1439_ngat) );
INVXL U_g3712 (.A(G3959GAT_1440_gat), .Y(G3959GAT_1440_ngat) );
INVXL U_g3713 (.A(G3955GAT_1441_gat), .Y(G3955GAT_1441_ngat) );
INVXL U_g3714 (.A(G3951GAT_1442_gat), .Y(G3951GAT_1442_ngat) );
INVXL U_g3715 (.A(G3947GAT_1443_gat), .Y(G3947GAT_1443_ngat) );
INVXL U_g3716 (.A(G3977GAT_1431_gat), .Y(G3977GAT_1431_ngat) );
INVXL U_g3717 (.A(G954GAT_150_gat), .Y(G954GAT_150_ngat) );
INVXL U_g3718 (.A(G1293GAT_37_gat), .Y(G1293GAT_37_ngat) );
INVXL U_g3719 (.A(G4049GAT_1444_gat), .Y(G4049GAT_1444_ngat) );
INVXL U_g3720 (.A(G4047GAT_1445_gat), .Y(G4047GAT_1445_ngat) );
INVXL U_g3721 (.A(G4048GAT_1455_gat), .Y(G4048GAT_1455_ngat) );
INVXL U_g3722 (.A(G4043GAT_1457_gat), .Y(G4043GAT_1457_ngat) );
INVXL U_g3723 (.A(G4038GAT_1447_gat), .Y(G4038GAT_1447_ngat) );
INVXL U_g3724 (.A(G4039GAT_1448_gat), .Y(G4039GAT_1448_ngat) );
INVXL U_g3725 (.A(G4034GAT_1449_gat), .Y(G4034GAT_1449_ngat) );
INVXL U_g3726 (.A(G4031GAT_1450_gat), .Y(G4031GAT_1450_ngat) );
INVXL U_g3727 (.A(G4028GAT_1451_gat), .Y(G4028GAT_1451_ngat) );
INVXL U_g3728 (.A(G4026GAT_1452_gat), .Y(G4026GAT_1452_ngat) );
INVXL U_g3729 (.A(G4027GAT_1462_gat), .Y(G4027GAT_1462_ngat) );
INVXL U_g3730 (.A(G4022GAT_1464_gat), .Y(G4022GAT_1464_ngat) );
INVXL U_g3731 (.A(G4017GAT_1454_gat), .Y(G4017GAT_1454_ngat) );
INVXL U_g3732 (.A(G4018GAT_1465_gat), .Y(G4018GAT_1465_ngat) );
INVXL U_g3733 (.A(G4015GAT_1456_gat), .Y(G4015GAT_1456_ngat) );
INVXL U_g3734 (.A(G4016GAT_1466_gat), .Y(G4016GAT_1466_ngat) );
INVXL U_g3735 (.A(G4013GAT_1458_gat), .Y(G4013GAT_1458_ngat) );
INVXL U_g3736 (.A(G4014GAT_1467_gat), .Y(G4014GAT_1467_ngat) );
INVXL U_g3737 (.A(G4040GAT_1446_gat), .Y(G4040GAT_1446_ngat) );
INVXL U_g3738 (.A(G1149GAT_85_gat), .Y(G1149GAT_85_ngat) );
INVXL U_g3739 (.A(G4011GAT_1459_gat), .Y(G4011GAT_1459_ngat) );
INVXL U_g3740 (.A(G4012GAT_1468_gat), .Y(G4012GAT_1468_ngat) );
INVXL U_g3741 (.A(G4009GAT_1460_gat), .Y(G4009GAT_1460_ngat) );
INVXL U_g3742 (.A(G4010GAT_1469_gat), .Y(G4010GAT_1469_ngat) );
INVXL U_g3743 (.A(G4007GAT_1461_gat), .Y(G4007GAT_1461_ngat) );
INVXL U_g3744 (.A(G4008GAT_1470_gat), .Y(G4008GAT_1470_ngat) );
INVXL U_g3745 (.A(G4005GAT_1463_gat), .Y(G4005GAT_1463_ngat) );
INVXL U_g3746 (.A(G4006GAT_1471_gat), .Y(G4006GAT_1471_ngat) );
INVXL U_g3747 (.A(G4019GAT_1453_gat), .Y(G4019GAT_1453_ngat) );
INVXL U_g3748 (.A(G906GAT_166_gat), .Y(G906GAT_166_ngat) );
INVXL U_g3749 (.A(G4106GAT_1472_gat), .Y(G4106GAT_1472_ngat) );
INVXL U_g3750 (.A(G4103GAT_1473_gat), .Y(G4103GAT_1473_ngat) );
INVXL U_g3751 (.A(G4100GAT_1474_gat), .Y(G4100GAT_1474_ngat) );
INVXL U_g3752 (.A(G4098GAT_1475_gat), .Y(G4098GAT_1475_ngat) );
INVXL U_g3753 (.A(G4099GAT_1485_gat), .Y(G4099GAT_1485_ngat) );
INVXL U_g3754 (.A(G4094GAT_1487_gat), .Y(G4094GAT_1487_ngat) );
INVXL U_g3755 (.A(G4089GAT_1477_gat), .Y(G4089GAT_1477_ngat) );
INVXL U_g3756 (.A(G4090GAT_1478_gat), .Y(G4090GAT_1478_ngat) );
INVXL U_g3757 (.A(G4085GAT_1479_gat), .Y(G4085GAT_1479_ngat) );
INVXL U_g3758 (.A(G4082GAT_1480_gat), .Y(G4082GAT_1480_ngat) );
INVXL U_g3759 (.A(G4079GAT_1481_gat), .Y(G4079GAT_1481_ngat) );
INVXL U_g3760 (.A(G4077GAT_1482_gat), .Y(G4077GAT_1482_ngat) );
INVXL U_g3761 (.A(G4078GAT_1492_gat), .Y(G4078GAT_1492_ngat) );
INVXL U_g3762 (.A(G4073GAT_1493_gat), .Y(G4073GAT_1493_ngat) );
INVXL U_g3763 (.A(G4091GAT_1476_gat), .Y(G4091GAT_1476_ngat) );
INVXL U_g3764 (.A(G1101GAT_101_gat), .Y(G1101GAT_101_ngat) );
INVXL U_g3765 (.A(G4070GAT_1483_gat), .Y(G4070GAT_1483_ngat) );
INVXL U_g3766 (.A(G858GAT_182_gat), .Y(G858GAT_182_ngat) );
INVXL U_g3767 (.A(G4067GAT_1484_gat), .Y(G4067GAT_1484_ngat) );
INVXL U_g3768 (.A(G810GAT_198_gat), .Y(G810GAT_198_ngat) );
INVXL U_g3769 (.A(G4064GAT_1486_gat), .Y(G4064GAT_1486_ngat) );
INVXL U_g3770 (.A(G762GAT_214_gat), .Y(G762GAT_214_ngat) );
INVXL U_g3771 (.A(G4061GAT_1488_gat), .Y(G4061GAT_1488_ngat) );
INVXL U_g3772 (.A(G714GAT_230_gat), .Y(G714GAT_230_ngat) );
INVXL U_g3773 (.A(G4058GAT_1489_gat), .Y(G4058GAT_1489_ngat) );
INVXL U_g3774 (.A(G666GAT_246_gat), .Y(G666GAT_246_ngat) );
INVXL U_g3775 (.A(G4055GAT_1490_gat), .Y(G4055GAT_1490_ngat) );
INVXL U_g3776 (.A(G618GAT_262_gat), .Y(G618GAT_262_ngat) );
INVXL U_g3777 (.A(G4052GAT_1491_gat), .Y(G4052GAT_1491_ngat) );
INVXL U_g3778 (.A(G570GAT_278_gat), .Y(G570GAT_278_ngat) );
INVXL U_g3779 (.A(G4171GAT_1494_gat), .Y(G4171GAT_1494_ngat) );
INVXL U_g3780 (.A(G4172GAT_1495_gat), .Y(G4172GAT_1495_ngat) );
INVXL U_g3781 (.A(G4167GAT_1496_gat), .Y(G4167GAT_1496_ngat) );
INVXL U_g3782 (.A(G4164GAT_1497_gat), .Y(G4164GAT_1497_ngat) );
INVXL U_g3783 (.A(G4161GAT_1498_gat), .Y(G4161GAT_1498_ngat) );
INVXL U_g3784 (.A(G4159GAT_1499_gat), .Y(G4159GAT_1499_ngat) );
INVXL U_g3785 (.A(G4160GAT_1507_gat), .Y(G4160GAT_1507_ngat) );
INVXL U_g3786 (.A(G4155GAT_1508_gat), .Y(G4155GAT_1508_ngat) );
INVXL U_g3787 (.A(G4150GAT_1501_gat), .Y(G4150GAT_1501_ngat) );
INVXL U_g3788 (.A(G4151GAT_1502_gat), .Y(G4151GAT_1502_ngat) );
INVXL U_g3789 (.A(G4146GAT_1503_gat), .Y(G4146GAT_1503_ngat) );
INVXL U_g3790 (.A(G4143GAT_1504_gat), .Y(G4143GAT_1504_ngat) );
INVXL U_g3791 (.A(G4140GAT_1505_gat), .Y(G4140GAT_1505_ngat) );
INVXL U_g3792 (.A(G4138GAT_1506_gat), .Y(G4138GAT_1506_ngat) );
INVXL U_g3793 (.A(G4139GAT_1509_gat), .Y(G4139GAT_1509_ngat) );
INVXL U_g3794 (.A(G4134GAT_1510_gat), .Y(G4134GAT_1510_ngat) );
INVXL U_g3795 (.A(G4130GAT_1511_gat), .Y(G4130GAT_1511_ngat) );
INVXL U_g3796 (.A(G4126GAT_1512_gat), .Y(G4126GAT_1512_ngat) );
INVXL U_g3797 (.A(G4122GAT_1513_gat), .Y(G4122GAT_1513_ngat) );
INVXL U_g3798 (.A(G4118GAT_1514_gat), .Y(G4118GAT_1514_ngat) );
INVXL U_g3799 (.A(G4152GAT_1500_gat), .Y(G4152GAT_1500_ngat) );
INVXL U_g3800 (.A(G1053GAT_117_gat), .Y(G1053GAT_117_ngat) );
INVXL U_g3801 (.A(G4114GAT_1515_gat), .Y(G4114GAT_1515_ngat) );
INVXL U_g3802 (.A(G4110GAT_1516_gat), .Y(G4110GAT_1516_ngat) );
INVXL U_g3803 (.A(G4236GAT_1518_gat), .Y(G4236GAT_1518_ngat) );
INVXL U_g3804 (.A(G4237GAT_1519_gat), .Y(G4237GAT_1519_ngat) );
INVXL U_g3805 (.A(G4232GAT_1520_gat), .Y(G4232GAT_1520_ngat) );
INVXL U_g3806 (.A(G4229GAT_1521_gat), .Y(G4229GAT_1521_ngat) );
INVXL U_g3807 (.A(G4226GAT_1522_gat), .Y(G4226GAT_1522_ngat) );
INVXL U_g3808 (.A(G4224GAT_1523_gat), .Y(G4224GAT_1523_ngat) );
INVXL U_g3809 (.A(G4225GAT_1533_gat), .Y(G4225GAT_1533_ngat) );
INVXL U_g3810 (.A(G4220GAT_1535_gat), .Y(G4220GAT_1535_ngat) );
INVXL U_g3811 (.A(G4215GAT_1525_gat), .Y(G4215GAT_1525_ngat) );
INVXL U_g3812 (.A(G4216GAT_1526_gat), .Y(G4216GAT_1526_ngat) );
INVXL U_g3813 (.A(G4211GAT_1527_gat), .Y(G4211GAT_1527_ngat) );
INVXL U_g3814 (.A(G4208GAT_1528_gat), .Y(G4208GAT_1528_ngat) );
INVXL U_g3815 (.A(G4205GAT_1538_gat), .Y(G4205GAT_1538_ngat) );
INVXL U_g3816 (.A(G4203GAT_1529_gat), .Y(G4203GAT_1529_ngat) );
INVXL U_g3817 (.A(G4204GAT_1539_gat), .Y(G4204GAT_1539_ngat) );
INVXL U_g3818 (.A(G4238GAT_1517_gat), .Y(G4238GAT_1517_ngat) );
INVXL U_g3819 (.A(G1248GAT_52_gat), .Y(G1248GAT_52_ngat) );
INVXL U_g3820 (.A(G4198GAT_1530_gat), .Y(G4198GAT_1530_ngat) );
INVXL U_g3821 (.A(G4199GAT_1541_gat), .Y(G4199GAT_1541_ngat) );
INVXL U_g3822 (.A(G4193GAT_1531_gat), .Y(G4193GAT_1531_ngat) );
INVXL U_g3823 (.A(G4194GAT_1543_gat), .Y(G4194GAT_1543_ngat) );
INVXL U_g3824 (.A(G4188GAT_1532_gat), .Y(G4188GAT_1532_ngat) );
INVXL U_g3825 (.A(G4189GAT_1545_gat), .Y(G4189GAT_1545_ngat) );
INVXL U_g3826 (.A(G4183GAT_1534_gat), .Y(G4183GAT_1534_ngat) );
INVXL U_g3827 (.A(G4184GAT_1547_gat), .Y(G4184GAT_1547_ngat) );
INVXL U_g3828 (.A(G4178GAT_1536_gat), .Y(G4178GAT_1536_ngat) );
INVXL U_g3829 (.A(G4179GAT_1549_gat), .Y(G4179GAT_1549_ngat) );
INVXL U_g3830 (.A(G4217GAT_1524_gat), .Y(G4217GAT_1524_ngat) );
INVXL U_g3831 (.A(G1005GAT_133_gat), .Y(G1005GAT_133_ngat) );
INVXL U_g3832 (.A(G4173GAT_1537_gat), .Y(G4173GAT_1537_ngat) );
INVXL U_g3833 (.A(G4174GAT_1551_gat), .Y(G4174GAT_1551_ngat) );
INVXL U_g3834 (.A(G4290GAT_1564_gat), .Y(G4290GAT_1564_ngat) );
INVXL U_g3835 (.A(G4285GAT_1553_gat), .Y(G4285GAT_1553_ngat) );
INVXL U_g3836 (.A(G4286GAT_1554_gat), .Y(G4286GAT_1554_ngat) );
INVXL U_g3837 (.A(G4281GAT_1555_gat), .Y(G4281GAT_1555_ngat) );
INVXL U_g3838 (.A(G4278GAT_1556_gat), .Y(G4278GAT_1556_ngat) );
INVXL U_g3839 (.A(G4275GAT_1557_gat), .Y(G4275GAT_1557_ngat) );
INVXL U_g3840 (.A(G4273GAT_1558_gat), .Y(G4273GAT_1558_ngat) );
INVXL U_g3841 (.A(G4274GAT_1569_gat), .Y(G4274GAT_1569_ngat) );
INVXL U_g3842 (.A(G4269GAT_1571_gat), .Y(G4269GAT_1571_ngat) );
INVXL U_g3843 (.A(G4264GAT_1560_gat), .Y(G4264GAT_1560_ngat) );
INVXL U_g3844 (.A(G4265GAT_1561_gat), .Y(G4265GAT_1561_ngat) );
INVXL U_g3845 (.A(G4260GAT_1562_gat), .Y(G4260GAT_1562_ngat) );
INVXL U_g3846 (.A(G4287GAT_1552_gat), .Y(G4287GAT_1552_ngat) );
INVXL U_g3847 (.A(G1200GAT_68_gat), .Y(G1200GAT_68_ngat) );
INVXL U_g3848 (.A(G4266GAT_1559_gat), .Y(G4266GAT_1559_ngat) );
INVXL U_g3849 (.A(G957GAT_149_gat), .Y(G957GAT_149_ngat) );
INVXL U_g3850 (.A(G4257GAT_1563_gat), .Y(G4257GAT_1563_ngat) );
INVXL U_g3851 (.A(G4200GAT_1540_gat), .Y(G4200GAT_1540_ngat) );
INVXL U_g3852 (.A(G4254GAT_1565_gat), .Y(G4254GAT_1565_ngat) );
INVXL U_g3853 (.A(G4195GAT_1542_gat), .Y(G4195GAT_1542_ngat) );
INVXL U_g3854 (.A(G4251GAT_1566_gat), .Y(G4251GAT_1566_ngat) );
INVXL U_g3855 (.A(G4190GAT_1544_gat), .Y(G4190GAT_1544_ngat) );
INVXL U_g3856 (.A(G4248GAT_1567_gat), .Y(G4248GAT_1567_ngat) );
INVXL U_g3857 (.A(G4185GAT_1546_gat), .Y(G4185GAT_1546_ngat) );
INVXL U_g3858 (.A(G4245GAT_1568_gat), .Y(G4245GAT_1568_ngat) );
INVXL U_g3859 (.A(G4180GAT_1548_gat), .Y(G4180GAT_1548_ngat) );
INVXL U_g3860 (.A(G4242GAT_1570_gat), .Y(G4242GAT_1570_ngat) );
INVXL U_g3861 (.A(G4175GAT_1550_gat), .Y(G4175GAT_1550_ngat) );
INVXL U_g3862 (.A(G1296GAT_36_gat), .Y(G1296GAT_36_ngat) );
INVXL U_g3863 (.A(G4350GAT_1573_gat), .Y(G4350GAT_1573_ngat) );
INVXL U_g3864 (.A(G4348GAT_1574_gat), .Y(G4348GAT_1574_ngat) );
INVXL U_g3865 (.A(G4349GAT_1584_gat), .Y(G4349GAT_1584_ngat) );
INVXL U_g3866 (.A(G4344GAT_1585_gat), .Y(G4344GAT_1585_ngat) );
INVXL U_g3867 (.A(G4339GAT_1576_gat), .Y(G4339GAT_1576_ngat) );
INVXL U_g3868 (.A(G4340GAT_1577_gat), .Y(G4340GAT_1577_ngat) );
INVXL U_g3869 (.A(G4335GAT_1578_gat), .Y(G4335GAT_1578_ngat) );
INVXL U_g3870 (.A(G4332GAT_1579_gat), .Y(G4332GAT_1579_ngat) );
INVXL U_g3871 (.A(G4329GAT_1580_gat), .Y(G4329GAT_1580_ngat) );
INVXL U_g3872 (.A(G4327GAT_1581_gat), .Y(G4327GAT_1581_ngat) );
INVXL U_g3873 (.A(G4328GAT_1586_gat), .Y(G4328GAT_1586_ngat) );
INVXL U_g3874 (.A(G4323GAT_1587_gat), .Y(G4323GAT_1587_ngat) );
INVXL U_g3875 (.A(G4318GAT_1583_gat), .Y(G4318GAT_1583_ngat) );
INVXL U_g3876 (.A(G4319GAT_1588_gat), .Y(G4319GAT_1588_ngat) );
INVXL U_g3877 (.A(G4314GAT_1589_gat), .Y(G4314GAT_1589_ngat) );
INVXL U_g3878 (.A(G4310GAT_1590_gat), .Y(G4310GAT_1590_ngat) );
INVXL U_g3879 (.A(G4306GAT_1591_gat), .Y(G4306GAT_1591_ngat) );
INVXL U_g3880 (.A(G4341GAT_1575_gat), .Y(G4341GAT_1575_ngat) );
INVXL U_g3881 (.A(G1152GAT_84_gat), .Y(G1152GAT_84_ngat) );
INVXL U_g3882 (.A(G4302GAT_1592_gat), .Y(G4302GAT_1592_ngat) );
INVXL U_g3883 (.A(G4298GAT_1593_gat), .Y(G4298GAT_1593_ngat) );
INVXL U_g3884 (.A(G4294GAT_1594_gat), .Y(G4294GAT_1594_ngat) );
INVXL U_g3885 (.A(G4320GAT_1582_gat), .Y(G4320GAT_1582_ngat) );
INVXL U_g3886 (.A(G909GAT_165_gat), .Y(G909GAT_165_ngat) );
INVXL U_g3887 (.A(G4401GAT_1595_gat), .Y(G4401GAT_1595_ngat) );
INVXL U_g3888 (.A(G4398GAT_1596_gat), .Y(G4398GAT_1596_ngat) );
INVXL U_g3889 (.A(G4395GAT_1597_gat), .Y(G4395GAT_1597_ngat) );
INVXL U_g3890 (.A(G4393GAT_1598_gat), .Y(G4393GAT_1598_ngat) );
INVXL U_g3891 (.A(G4394GAT_1609_gat), .Y(G4394GAT_1609_ngat) );
INVXL U_g3892 (.A(G4389GAT_1611_gat), .Y(G4389GAT_1611_ngat) );
INVXL U_g3893 (.A(G4384GAT_1600_gat), .Y(G4384GAT_1600_ngat) );
INVXL U_g3894 (.A(G4385GAT_1601_gat), .Y(G4385GAT_1601_ngat) );
INVXL U_g3895 (.A(G4380GAT_1602_gat), .Y(G4380GAT_1602_ngat) );
INVXL U_g3896 (.A(G4377GAT_1603_gat), .Y(G4377GAT_1603_ngat) );
INVXL U_g3897 (.A(G4374GAT_1604_gat), .Y(G4374GAT_1604_ngat) );
INVXL U_g3898 (.A(G4372GAT_1605_gat), .Y(G4372GAT_1605_ngat) );
INVXL U_g3899 (.A(G4373GAT_1615_gat), .Y(G4373GAT_1615_ngat) );
INVXL U_g3900 (.A(G4368GAT_1616_gat), .Y(G4368GAT_1616_ngat) );
INVXL U_g3901 (.A(G4363GAT_1607_gat), .Y(G4363GAT_1607_ngat) );
INVXL U_g3902 (.A(G4364GAT_1617_gat), .Y(G4364GAT_1617_ngat) );
INVXL U_g3903 (.A(G4361GAT_1608_gat), .Y(G4361GAT_1608_ngat) );
INVXL U_g3904 (.A(G4362GAT_1618_gat), .Y(G4362GAT_1618_ngat) );
INVXL U_g3905 (.A(G4359GAT_1610_gat), .Y(G4359GAT_1610_ngat) );
INVXL U_g3906 (.A(G4360GAT_1619_gat), .Y(G4360GAT_1619_ngat) );
INVXL U_g3907 (.A(G4357GAT_1612_gat), .Y(G4357GAT_1612_ngat) );
INVXL U_g3908 (.A(G4358GAT_1620_gat), .Y(G4358GAT_1620_ngat) );
INVXL U_g3909 (.A(G4386GAT_1599_gat), .Y(G4386GAT_1599_ngat) );
INVXL U_g3910 (.A(G1104GAT_100_gat), .Y(G1104GAT_100_ngat) );
INVXL U_g3911 (.A(G4355GAT_1613_gat), .Y(G4355GAT_1613_ngat) );
INVXL U_g3912 (.A(G4356GAT_1621_gat), .Y(G4356GAT_1621_ngat) );
INVXL U_g3913 (.A(G4353GAT_1614_gat), .Y(G4353GAT_1614_ngat) );
INVXL U_g3914 (.A(G4354GAT_1622_gat), .Y(G4354GAT_1622_ngat) );
INVXL U_g3915 (.A(G4365GAT_1606_gat), .Y(G4365GAT_1606_ngat) );
INVXL U_g3916 (.A(G861GAT_181_gat), .Y(G861GAT_181_ngat) );
INVXL U_g3917 (.A(G4460GAT_1623_gat), .Y(G4460GAT_1623_ngat) );
INVXL U_g3918 (.A(G4461GAT_1624_gat), .Y(G4461GAT_1624_ngat) );
INVXL U_g3919 (.A(G4456GAT_1625_gat), .Y(G4456GAT_1625_ngat) );
INVXL U_g3920 (.A(G4453GAT_1626_gat), .Y(G4453GAT_1626_ngat) );
INVXL U_g3921 (.A(G4450GAT_1627_gat), .Y(G4450GAT_1627_ngat) );
INVXL U_g3922 (.A(G4448GAT_1628_gat), .Y(G4448GAT_1628_ngat) );
INVXL U_g3923 (.A(G4449GAT_1639_gat), .Y(G4449GAT_1639_ngat) );
INVXL U_g3924 (.A(G4444GAT_1641_gat), .Y(G4444GAT_1641_ngat) );
INVXL U_g3925 (.A(G4439GAT_1630_gat), .Y(G4439GAT_1630_ngat) );
INVXL U_g3926 (.A(G4440GAT_1631_gat), .Y(G4440GAT_1631_ngat) );
INVXL U_g3927 (.A(G4435GAT_1632_gat), .Y(G4435GAT_1632_ngat) );
INVXL U_g3928 (.A(G4432GAT_1633_gat), .Y(G4432GAT_1633_ngat) );
INVXL U_g3929 (.A(G4429GAT_1634_gat), .Y(G4429GAT_1634_ngat) );
INVXL U_g3930 (.A(G4427GAT_1635_gat), .Y(G4427GAT_1635_ngat) );
INVXL U_g3931 (.A(G4428GAT_1644_gat), .Y(G4428GAT_1644_ngat) );
INVXL U_g3932 (.A(G4423GAT_1645_gat), .Y(G4423GAT_1645_ngat) );
INVXL U_g3933 (.A(G4441GAT_1629_gat), .Y(G4441GAT_1629_ngat) );
INVXL U_g3934 (.A(G1056GAT_116_gat), .Y(G1056GAT_116_ngat) );
INVXL U_g3935 (.A(G4420GAT_1636_gat), .Y(G4420GAT_1636_ngat) );
INVXL U_g3936 (.A(G813GAT_197_gat), .Y(G813GAT_197_ngat) );
INVXL U_g3937 (.A(G4417GAT_1637_gat), .Y(G4417GAT_1637_ngat) );
INVXL U_g3938 (.A(G765GAT_213_gat), .Y(G765GAT_213_ngat) );
INVXL U_g3939 (.A(G4414GAT_1638_gat), .Y(G4414GAT_1638_ngat) );
INVXL U_g3940 (.A(G717GAT_229_gat), .Y(G717GAT_229_ngat) );
INVXL U_g3941 (.A(G4411GAT_1640_gat), .Y(G4411GAT_1640_ngat) );
INVXL U_g3942 (.A(G669GAT_245_gat), .Y(G669GAT_245_ngat) );
INVXL U_g3943 (.A(G4408GAT_1642_gat), .Y(G4408GAT_1642_ngat) );
INVXL U_g3944 (.A(G621GAT_261_gat), .Y(G621GAT_261_ngat) );
INVXL U_g3945 (.A(G4405GAT_1643_gat), .Y(G4405GAT_1643_ngat) );
INVXL U_g3946 (.A(G573GAT_277_gat), .Y(G573GAT_277_ngat) );
INVXL U_g3947 (.A(G4519GAT_1647_gat), .Y(G4519GAT_1647_ngat) );
INVXL U_g3948 (.A(G4520GAT_1648_gat), .Y(G4520GAT_1648_ngat) );
INVXL U_g3949 (.A(G4515GAT_1649_gat), .Y(G4515GAT_1649_ngat) );
INVXL U_g3950 (.A(G4512GAT_1650_gat), .Y(G4512GAT_1650_ngat) );
INVXL U_g3951 (.A(G4509GAT_1651_gat), .Y(G4509GAT_1651_ngat) );
INVXL U_g3952 (.A(G4507GAT_1652_gat), .Y(G4507GAT_1652_ngat) );
INVXL U_g3953 (.A(G4508GAT_1660_gat), .Y(G4508GAT_1660_ngat) );
INVXL U_g3954 (.A(G4503GAT_1661_gat), .Y(G4503GAT_1661_ngat) );
INVXL U_g3955 (.A(G4498GAT_1654_gat), .Y(G4498GAT_1654_ngat) );
INVXL U_g3956 (.A(G4499GAT_1655_gat), .Y(G4499GAT_1655_ngat) );
INVXL U_g3957 (.A(G4494GAT_1656_gat), .Y(G4494GAT_1656_ngat) );
INVXL U_g3958 (.A(G4491GAT_1657_gat), .Y(G4491GAT_1657_ngat) );
INVXL U_g3959 (.A(G4488GAT_1658_gat), .Y(G4488GAT_1658_ngat) );
INVXL U_g3960 (.A(G4486GAT_1659_gat), .Y(G4486GAT_1659_ngat) );
INVXL U_g3961 (.A(G4487GAT_1662_gat), .Y(G4487GAT_1662_ngat) );
INVXL U_g3962 (.A(G4482GAT_1663_gat), .Y(G4482GAT_1663_ngat) );
INVXL U_g3963 (.A(G4521GAT_1646_gat), .Y(G4521GAT_1646_ngat) );
INVXL U_g3964 (.A(G1251GAT_51_gat), .Y(G1251GAT_51_ngat) );
INVXL U_g3965 (.A(G4478GAT_1664_gat), .Y(G4478GAT_1664_ngat) );
INVXL U_g3966 (.A(G4474GAT_1665_gat), .Y(G4474GAT_1665_ngat) );
INVXL U_g3967 (.A(G4470GAT_1666_gat), .Y(G4470GAT_1666_ngat) );
INVXL U_g3968 (.A(G4466GAT_1667_gat), .Y(G4466GAT_1667_ngat) );
INVXL U_g3969 (.A(G4462GAT_1668_gat), .Y(G4462GAT_1668_ngat) );
INVXL U_g3970 (.A(G4500GAT_1653_gat), .Y(G4500GAT_1653_ngat) );
INVXL U_g3971 (.A(G1008GAT_132_gat), .Y(G1008GAT_132_ngat) );
INVXL U_g3972 (.A(G4587GAT_1682_gat), .Y(G4587GAT_1682_ngat) );
INVXL U_g3973 (.A(G4582GAT_1670_gat), .Y(G4582GAT_1670_ngat) );
INVXL U_g3974 (.A(G4583GAT_1671_gat), .Y(G4583GAT_1671_ngat) );
INVXL U_g3975 (.A(G4578GAT_1672_gat), .Y(G4578GAT_1672_ngat) );
INVXL U_g3976 (.A(G4575GAT_1673_gat), .Y(G4575GAT_1673_ngat) );
INVXL U_g3977 (.A(G4572GAT_1674_gat), .Y(G4572GAT_1674_ngat) );
INVXL U_g3978 (.A(G4570GAT_1675_gat), .Y(G4570GAT_1675_ngat) );
INVXL U_g3979 (.A(G4571GAT_1687_gat), .Y(G4571GAT_1687_ngat) );
INVXL U_g3980 (.A(G4566GAT_1689_gat), .Y(G4566GAT_1689_ngat) );
INVXL U_g3981 (.A(G4561GAT_1677_gat), .Y(G4561GAT_1677_ngat) );
INVXL U_g3982 (.A(G4562GAT_1678_gat), .Y(G4562GAT_1678_ngat) );
INVXL U_g3983 (.A(G4557GAT_1679_gat), .Y(G4557GAT_1679_ngat) );
INVXL U_g3984 (.A(G4554GAT_1680_gat), .Y(G4554GAT_1680_ngat) );
INVXL U_g3985 (.A(G4551GAT_1690_gat), .Y(G4551GAT_1690_ngat) );
INVXL U_g3986 (.A(G4549GAT_1681_gat), .Y(G4549GAT_1681_ngat) );
INVXL U_g3987 (.A(G4550GAT_1691_gat), .Y(G4550GAT_1691_ngat) );
INVXL U_g3988 (.A(G4544GAT_1683_gat), .Y(G4544GAT_1683_ngat) );
INVXL U_g3989 (.A(G4545GAT_1693_gat), .Y(G4545GAT_1693_ngat) );
INVXL U_g3990 (.A(G4584GAT_1669_gat), .Y(G4584GAT_1669_ngat) );
INVXL U_g3991 (.A(G1203GAT_67_gat), .Y(G1203GAT_67_ngat) );
INVXL U_g3992 (.A(G4539GAT_1684_gat), .Y(G4539GAT_1684_ngat) );
INVXL U_g3993 (.A(G4540GAT_1695_gat), .Y(G4540GAT_1695_ngat) );
INVXL U_g3994 (.A(G4534GAT_1685_gat), .Y(G4534GAT_1685_ngat) );
INVXL U_g3995 (.A(G4535GAT_1697_gat), .Y(G4535GAT_1697_ngat) );
INVXL U_g3996 (.A(G4529GAT_1686_gat), .Y(G4529GAT_1686_ngat) );
INVXL U_g3997 (.A(G4530GAT_1699_gat), .Y(G4530GAT_1699_ngat) );
INVXL U_g3998 (.A(G4524GAT_1688_gat), .Y(G4524GAT_1688_ngat) );
INVXL U_g3999 (.A(G4525GAT_1701_gat), .Y(G4525GAT_1701_ngat) );
INVXL U_g4000 (.A(G4563GAT_1676_gat), .Y(G4563GAT_1676_ngat) );
INVXL U_g4001 (.A(G960GAT_148_gat), .Y(G960GAT_148_ngat) );
INVXL U_g4002 (.A(G1299GAT_35_gat), .Y(G1299GAT_35_ngat) );
INVXL U_g4003 (.A(G4643GAT_1702_gat), .Y(G4643GAT_1702_ngat) );
INVXL U_g4004 (.A(G4641GAT_1703_gat), .Y(G4641GAT_1703_ngat) );
INVXL U_g4005 (.A(G4642GAT_1716_gat), .Y(G4642GAT_1716_ngat) );
INVXL U_g4006 (.A(G4637GAT_1718_gat), .Y(G4637GAT_1718_ngat) );
INVXL U_g4007 (.A(G4632GAT_1705_gat), .Y(G4632GAT_1705_ngat) );
INVXL U_g4008 (.A(G4633GAT_1706_gat), .Y(G4633GAT_1706_ngat) );
INVXL U_g4009 (.A(G4628GAT_1707_gat), .Y(G4628GAT_1707_ngat) );
INVXL U_g4010 (.A(G4625GAT_1708_gat), .Y(G4625GAT_1708_ngat) );
INVXL U_g4011 (.A(G4622GAT_1709_gat), .Y(G4622GAT_1709_ngat) );
INVXL U_g4012 (.A(G4620GAT_1710_gat), .Y(G4620GAT_1710_ngat) );
INVXL U_g4013 (.A(G4621GAT_1723_gat), .Y(G4621GAT_1723_ngat) );
INVXL U_g4014 (.A(G4616GAT_1724_gat), .Y(G4616GAT_1724_ngat) );
INVXL U_g4015 (.A(G4611GAT_1712_gat), .Y(G4611GAT_1712_ngat) );
INVXL U_g4016 (.A(G4612GAT_1713_gat), .Y(G4612GAT_1713_ngat) );
INVXL U_g4017 (.A(G4607GAT_1714_gat), .Y(G4607GAT_1714_ngat) );
INVXL U_g4018 (.A(G4634GAT_1704_gat), .Y(G4634GAT_1704_ngat) );
INVXL U_g4019 (.A(G1155GAT_83_gat), .Y(G1155GAT_83_ngat) );
INVXL U_g4020 (.A(G4613GAT_1711_gat), .Y(G4613GAT_1711_ngat) );
INVXL U_g4021 (.A(G912GAT_164_gat), .Y(G912GAT_164_ngat) );
INVXL U_g4022 (.A(G4604GAT_1715_gat), .Y(G4604GAT_1715_ngat) );
INVXL U_g4023 (.A(G4546GAT_1692_gat), .Y(G4546GAT_1692_ngat) );
INVXL U_g4024 (.A(G4601GAT_1717_gat), .Y(G4601GAT_1717_ngat) );
INVXL U_g4025 (.A(G4541GAT_1694_gat), .Y(G4541GAT_1694_ngat) );
INVXL U_g4026 (.A(G4598GAT_1719_gat), .Y(G4598GAT_1719_ngat) );
INVXL U_g4027 (.A(G4536GAT_1696_gat), .Y(G4536GAT_1696_ngat) );
INVXL U_g4028 (.A(G4595GAT_1720_gat), .Y(G4595GAT_1720_ngat) );
INVXL U_g4029 (.A(G4531GAT_1698_gat), .Y(G4531GAT_1698_ngat) );
INVXL U_g4030 (.A(G4592GAT_1721_gat), .Y(G4592GAT_1721_ngat) );
INVXL U_g4031 (.A(G4526GAT_1700_gat), .Y(G4526GAT_1700_ngat) );
INVXL U_g4032 (.A(G4704GAT_1725_gat), .Y(G4704GAT_1725_ngat) );
INVXL U_g4033 (.A(G4701GAT_1726_gat), .Y(G4701GAT_1726_ngat) );
INVXL U_g4034 (.A(G4698GAT_1727_gat), .Y(G4698GAT_1727_ngat) );
INVXL U_g4035 (.A(G4696GAT_1728_gat), .Y(G4696GAT_1728_ngat) );
INVXL U_g4036 (.A(G4697GAT_1738_gat), .Y(G4697GAT_1738_ngat) );
INVXL U_g4037 (.A(G4692GAT_1739_gat), .Y(G4692GAT_1739_ngat) );
INVXL U_g4038 (.A(G4687GAT_1730_gat), .Y(G4687GAT_1730_ngat) );
INVXL U_g4039 (.A(G4688GAT_1731_gat), .Y(G4688GAT_1731_ngat) );
INVXL U_g4040 (.A(G4683GAT_1732_gat), .Y(G4683GAT_1732_ngat) );
INVXL U_g4041 (.A(G4680GAT_1733_gat), .Y(G4680GAT_1733_ngat) );
INVXL U_g4042 (.A(G4677GAT_1734_gat), .Y(G4677GAT_1734_ngat) );
INVXL U_g4043 (.A(G4675GAT_1735_gat), .Y(G4675GAT_1735_ngat) );
INVXL U_g4044 (.A(G4676GAT_1740_gat), .Y(G4676GAT_1740_ngat) );
INVXL U_g4045 (.A(G4671GAT_1741_gat), .Y(G4671GAT_1741_ngat) );
INVXL U_g4046 (.A(G4666GAT_1737_gat), .Y(G4666GAT_1737_ngat) );
INVXL U_g4047 (.A(G4667GAT_1742_gat), .Y(G4667GAT_1742_ngat) );
INVXL U_g4048 (.A(G4662GAT_1743_gat), .Y(G4662GAT_1743_ngat) );
INVXL U_g4049 (.A(G4658GAT_1744_gat), .Y(G4658GAT_1744_ngat) );
INVXL U_g4050 (.A(G4654GAT_1745_gat), .Y(G4654GAT_1745_ngat) );
INVXL U_g4051 (.A(G4650GAT_1746_gat), .Y(G4650GAT_1746_ngat) );
INVXL U_g4052 (.A(G4689GAT_1729_gat), .Y(G4689GAT_1729_ngat) );
INVXL U_g4053 (.A(G1107GAT_99_gat), .Y(G1107GAT_99_ngat) );
INVXL U_g4054 (.A(G4646GAT_1747_gat), .Y(G4646GAT_1747_ngat) );
INVXL U_g4055 (.A(G4668GAT_1736_gat), .Y(G4668GAT_1736_ngat) );
INVXL U_g4056 (.A(G864GAT_180_gat), .Y(G864GAT_180_ngat) );
INVXL U_g4057 (.A(G4758GAT_1748_gat), .Y(G4758GAT_1748_ngat) );
INVXL U_g4058 (.A(G4759GAT_1749_gat), .Y(G4759GAT_1749_ngat) );
INVXL U_g4059 (.A(G4754GAT_1750_gat), .Y(G4754GAT_1750_ngat) );
INVXL U_g4060 (.A(G4751GAT_1751_gat), .Y(G4751GAT_1751_ngat) );
INVXL U_g4061 (.A(G4748GAT_1752_gat), .Y(G4748GAT_1752_ngat) );
INVXL U_g4062 (.A(G4746GAT_1753_gat), .Y(G4746GAT_1753_ngat) );
INVXL U_g4063 (.A(G4747GAT_1765_gat), .Y(G4747GAT_1765_ngat) );
INVXL U_g4064 (.A(G4742GAT_1767_gat), .Y(G4742GAT_1767_ngat) );
INVXL U_g4065 (.A(G4737GAT_1755_gat), .Y(G4737GAT_1755_ngat) );
INVXL U_g4066 (.A(G4738GAT_1756_gat), .Y(G4738GAT_1756_ngat) );
INVXL U_g4067 (.A(G4733GAT_1757_gat), .Y(G4733GAT_1757_ngat) );
INVXL U_g4068 (.A(G4730GAT_1758_gat), .Y(G4730GAT_1758_ngat) );
INVXL U_g4069 (.A(G4727GAT_1759_gat), .Y(G4727GAT_1759_ngat) );
INVXL U_g4070 (.A(G4725GAT_1760_gat), .Y(G4725GAT_1760_ngat) );
INVXL U_g4071 (.A(G4726GAT_1769_gat), .Y(G4726GAT_1769_ngat) );
INVXL U_g4072 (.A(G4721GAT_1770_gat), .Y(G4721GAT_1770_ngat) );
INVXL U_g4073 (.A(G4716GAT_1762_gat), .Y(G4716GAT_1762_ngat) );
INVXL U_g4074 (.A(G4717GAT_1771_gat), .Y(G4717GAT_1771_ngat) );
INVXL U_g4075 (.A(G4714GAT_1763_gat), .Y(G4714GAT_1763_ngat) );
INVXL U_g4076 (.A(G4715GAT_1772_gat), .Y(G4715GAT_1772_ngat) );
INVXL U_g4077 (.A(G4712GAT_1764_gat), .Y(G4712GAT_1764_ngat) );
INVXL U_g4078 (.A(G4713GAT_1773_gat), .Y(G4713GAT_1773_ngat) );
INVXL U_g4079 (.A(G4710GAT_1766_gat), .Y(G4710GAT_1766_ngat) );
INVXL U_g4080 (.A(G4711GAT_1774_gat), .Y(G4711GAT_1774_ngat) );
INVXL U_g4081 (.A(G4708GAT_1768_gat), .Y(G4708GAT_1768_ngat) );
INVXL U_g4082 (.A(G4709GAT_1775_gat), .Y(G4709GAT_1775_ngat) );
INVXL U_g4083 (.A(G4739GAT_1754_gat), .Y(G4739GAT_1754_ngat) );
INVXL U_g4084 (.A(G1059GAT_115_gat), .Y(G1059GAT_115_ngat) );
INVXL U_g4085 (.A(G4718GAT_1761_gat), .Y(G4718GAT_1761_ngat) );
INVXL U_g4086 (.A(G816GAT_196_gat), .Y(G816GAT_196_ngat) );
INVXL U_g4087 (.A(G4812GAT_1777_gat), .Y(G4812GAT_1777_ngat) );
INVXL U_g4088 (.A(G4813GAT_1778_gat), .Y(G4813GAT_1778_ngat) );
INVXL U_g4089 (.A(G4808GAT_1779_gat), .Y(G4808GAT_1779_ngat) );
INVXL U_g4090 (.A(G4805GAT_1780_gat), .Y(G4805GAT_1780_ngat) );
INVXL U_g4091 (.A(G4802GAT_1781_gat), .Y(G4802GAT_1781_ngat) );
INVXL U_g4092 (.A(G4800GAT_1782_gat), .Y(G4800GAT_1782_ngat) );
INVXL U_g4093 (.A(G4801GAT_1794_gat), .Y(G4801GAT_1794_ngat) );
INVXL U_g4094 (.A(G4796GAT_1796_gat), .Y(G4796GAT_1796_ngat) );
INVXL U_g4095 (.A(G4791GAT_1784_gat), .Y(G4791GAT_1784_ngat) );
INVXL U_g4096 (.A(G4792GAT_1785_gat), .Y(G4792GAT_1785_ngat) );
INVXL U_g4097 (.A(G4787GAT_1786_gat), .Y(G4787GAT_1786_ngat) );
INVXL U_g4098 (.A(G4784GAT_1787_gat), .Y(G4784GAT_1787_ngat) );
INVXL U_g4099 (.A(G4781GAT_1788_gat), .Y(G4781GAT_1788_ngat) );
INVXL U_g4100 (.A(G4779GAT_1789_gat), .Y(G4779GAT_1789_ngat) );
INVXL U_g4101 (.A(G4780GAT_1797_gat), .Y(G4780GAT_1797_ngat) );
INVXL U_g4102 (.A(G4775GAT_1798_gat), .Y(G4775GAT_1798_ngat) );
INVXL U_g4103 (.A(G4814GAT_1776_gat), .Y(G4814GAT_1776_ngat) );
INVXL U_g4104 (.A(G1254GAT_50_gat), .Y(G1254GAT_50_ngat) );
INVXL U_g4105 (.A(G4793GAT_1783_gat), .Y(G4793GAT_1783_ngat) );
INVXL U_g4106 (.A(G1011GAT_131_gat), .Y(G1011GAT_131_ngat) );
INVXL U_g4107 (.A(G4772GAT_1790_gat), .Y(G4772GAT_1790_ngat) );
INVXL U_g4108 (.A(G768GAT_212_gat), .Y(G768GAT_212_ngat) );
INVXL U_g4109 (.A(G4769GAT_1791_gat), .Y(G4769GAT_1791_ngat) );
INVXL U_g4110 (.A(G720GAT_228_gat), .Y(G720GAT_228_ngat) );
INVXL U_g4111 (.A(G4766GAT_1792_gat), .Y(G4766GAT_1792_ngat) );
INVXL U_g4112 (.A(G672GAT_244_gat), .Y(G672GAT_244_ngat) );
INVXL U_g4113 (.A(G4763GAT_1793_gat), .Y(G4763GAT_1793_ngat) );
INVXL U_g4114 (.A(G624GAT_260_gat), .Y(G624GAT_260_ngat) );
INVXL U_g4115 (.A(G4760GAT_1795_gat), .Y(G4760GAT_1795_ngat) );
INVXL U_g4116 (.A(G576GAT_276_gat), .Y(G576GAT_276_ngat) );
INVXL U_g4117 (.A(G4875GAT_1813_gat), .Y(G4875GAT_1813_ngat) );
INVXL U_g4118 (.A(G4870GAT_1800_gat), .Y(G4870GAT_1800_ngat) );
INVXL U_g4119 (.A(G4871GAT_1801_gat), .Y(G4871GAT_1801_ngat) );
INVXL U_g4120 (.A(G4866GAT_1802_gat), .Y(G4866GAT_1802_ngat) );
INVXL U_g4121 (.A(G4863GAT_1803_gat), .Y(G4863GAT_1803_ngat) );
INVXL U_g4122 (.A(G4860GAT_1804_gat), .Y(G4860GAT_1804_ngat) );
INVXL U_g4123 (.A(G4858GAT_1805_gat), .Y(G4858GAT_1805_ngat) );
INVXL U_g4124 (.A(G4859GAT_1814_gat), .Y(G4859GAT_1814_ngat) );
INVXL U_g4125 (.A(G4854GAT_1815_gat), .Y(G4854GAT_1815_ngat) );
INVXL U_g4126 (.A(G4849GAT_1807_gat), .Y(G4849GAT_1807_ngat) );
INVXL U_g4127 (.A(G4850GAT_1808_gat), .Y(G4850GAT_1808_ngat) );
INVXL U_g4128 (.A(G4845GAT_1809_gat), .Y(G4845GAT_1809_ngat) );
INVXL U_g4129 (.A(G4842GAT_1810_gat), .Y(G4842GAT_1810_ngat) );
INVXL U_g4130 (.A(G4839GAT_1811_gat), .Y(G4839GAT_1811_ngat) );
INVXL U_g4131 (.A(G4837GAT_1812_gat), .Y(G4837GAT_1812_ngat) );
INVXL U_g4132 (.A(G4838GAT_1816_gat), .Y(G4838GAT_1816_ngat) );
INVXL U_g4133 (.A(G4833GAT_1817_gat), .Y(G4833GAT_1817_ngat) );
INVXL U_g4134 (.A(G4829GAT_1818_gat), .Y(G4829GAT_1818_ngat) );
INVXL U_g4135 (.A(G4872GAT_1799_gat), .Y(G4872GAT_1799_ngat) );
INVXL U_g4136 (.A(G1206GAT_66_gat), .Y(G1206GAT_66_ngat) );
INVXL U_g4137 (.A(G4825GAT_1819_gat), .Y(G4825GAT_1819_ngat) );
INVXL U_g4138 (.A(G4821GAT_1820_gat), .Y(G4821GAT_1820_ngat) );
INVXL U_g4139 (.A(G4817GAT_1821_gat), .Y(G4817GAT_1821_ngat) );
INVXL U_g4140 (.A(G4851GAT_1806_gat), .Y(G4851GAT_1806_ngat) );
INVXL U_g4141 (.A(G963GAT_147_gat), .Y(G963GAT_147_ngat) );
INVXL U_g4142 (.A(G1302GAT_34_gat), .Y(G1302GAT_34_ngat) );
INVXL U_g4143 (.A(G4943GAT_1822_gat), .Y(G4943GAT_1822_ngat) );
INVXL U_g4144 (.A(G4941GAT_1823_gat), .Y(G4941GAT_1823_ngat) );
INVXL U_g4145 (.A(G4942GAT_1837_gat), .Y(G4942GAT_1837_ngat) );
INVXL U_g4146 (.A(G4937GAT_1839_gat), .Y(G4937GAT_1839_ngat) );
INVXL U_g4147 (.A(G4932GAT_1825_gat), .Y(G4932GAT_1825_ngat) );
INVXL U_g4148 (.A(G4933GAT_1826_gat), .Y(G4933GAT_1826_ngat) );
INVXL U_g4149 (.A(G4928GAT_1827_gat), .Y(G4928GAT_1827_ngat) );
INVXL U_g4150 (.A(G4925GAT_1828_gat), .Y(G4925GAT_1828_ngat) );
INVXL U_g4151 (.A(G4922GAT_1829_gat), .Y(G4922GAT_1829_ngat) );
INVXL U_g4152 (.A(G4920GAT_1830_gat), .Y(G4920GAT_1830_ngat) );
INVXL U_g4153 (.A(G4921GAT_1843_gat), .Y(G4921GAT_1843_ngat) );
INVXL U_g4154 (.A(G4916GAT_1844_gat), .Y(G4916GAT_1844_ngat) );
INVXL U_g4155 (.A(G4911GAT_1832_gat), .Y(G4911GAT_1832_ngat) );
INVXL U_g4156 (.A(G4912GAT_1833_gat), .Y(G4912GAT_1833_ngat) );
INVXL U_g4157 (.A(G4907GAT_1834_gat), .Y(G4907GAT_1834_ngat) );
INVXL U_g4158 (.A(G4904GAT_1835_gat), .Y(G4904GAT_1835_ngat) );
INVXL U_g4159 (.A(G4901GAT_1845_gat), .Y(G4901GAT_1845_ngat) );
INVXL U_g4160 (.A(G4899GAT_1836_gat), .Y(G4899GAT_1836_ngat) );
INVXL U_g4161 (.A(G4900GAT_1846_gat), .Y(G4900GAT_1846_ngat) );
INVXL U_g4162 (.A(G4894GAT_1838_gat), .Y(G4894GAT_1838_ngat) );
INVXL U_g4163 (.A(G4895GAT_1848_gat), .Y(G4895GAT_1848_ngat) );
INVXL U_g4164 (.A(G4889GAT_1840_gat), .Y(G4889GAT_1840_ngat) );
INVXL U_g4165 (.A(G4890GAT_1850_gat), .Y(G4890GAT_1850_ngat) );
INVXL U_g4166 (.A(G4934GAT_1824_gat), .Y(G4934GAT_1824_ngat) );
INVXL U_g4167 (.A(G1158GAT_82_gat), .Y(G1158GAT_82_ngat) );
INVXL U_g4168 (.A(G4884GAT_1841_gat), .Y(G4884GAT_1841_ngat) );
INVXL U_g4169 (.A(G4885GAT_1852_gat), .Y(G4885GAT_1852_ngat) );
INVXL U_g4170 (.A(G4879GAT_1842_gat), .Y(G4879GAT_1842_ngat) );
INVXL U_g4171 (.A(G4880GAT_1854_gat), .Y(G4880GAT_1854_ngat) );
INVXL U_g4172 (.A(G4913GAT_1831_gat), .Y(G4913GAT_1831_ngat) );
INVXL U_g4173 (.A(G915GAT_163_gat), .Y(G915GAT_163_ngat) );
INVXL U_g4174 (.A(G5001GAT_1855_gat), .Y(G5001GAT_1855_ngat) );
INVXL U_g4175 (.A(G4998GAT_1856_gat), .Y(G4998GAT_1856_ngat) );
INVXL U_g4176 (.A(G4995GAT_1857_gat), .Y(G4995GAT_1857_ngat) );
INVXL U_g4177 (.A(G4993GAT_1858_gat), .Y(G4993GAT_1858_ngat) );
INVXL U_g4178 (.A(G4994GAT_1872_gat), .Y(G4994GAT_1872_ngat) );
INVXL U_g4179 (.A(G4989GAT_1874_gat), .Y(G4989GAT_1874_ngat) );
INVXL U_g4180 (.A(G4984GAT_1860_gat), .Y(G4984GAT_1860_ngat) );
INVXL U_g4181 (.A(G4985GAT_1861_gat), .Y(G4985GAT_1861_ngat) );
INVXL U_g4182 (.A(G4980GAT_1862_gat), .Y(G4980GAT_1862_ngat) );
INVXL U_g4183 (.A(G4977GAT_1863_gat), .Y(G4977GAT_1863_ngat) );
INVXL U_g4184 (.A(G4974GAT_1864_gat), .Y(G4974GAT_1864_ngat) );
INVXL U_g4185 (.A(G4972GAT_1865_gat), .Y(G4972GAT_1865_ngat) );
INVXL U_g4186 (.A(G4973GAT_1877_gat), .Y(G4973GAT_1877_ngat) );
INVXL U_g4187 (.A(G4968GAT_1878_gat), .Y(G4968GAT_1878_ngat) );
INVXL U_g4188 (.A(G4963GAT_1867_gat), .Y(G4963GAT_1867_ngat) );
INVXL U_g4189 (.A(G4964GAT_1868_gat), .Y(G4964GAT_1868_ngat) );
INVXL U_g4190 (.A(G4959GAT_1869_gat), .Y(G4959GAT_1869_ngat) );
INVXL U_g4191 (.A(G4986GAT_1859_gat), .Y(G4986GAT_1859_ngat) );
INVXL U_g4192 (.A(G1110GAT_98_gat), .Y(G1110GAT_98_ngat) );
INVXL U_g4193 (.A(G4965GAT_1866_gat), .Y(G4965GAT_1866_ngat) );
INVXL U_g4194 (.A(G867GAT_179_gat), .Y(G867GAT_179_ngat) );
INVXL U_g4195 (.A(G4956GAT_1870_gat), .Y(G4956GAT_1870_ngat) );
INVXL U_g4196 (.A(G4896GAT_1847_gat), .Y(G4896GAT_1847_ngat) );
INVXL U_g4197 (.A(G4953GAT_1871_gat), .Y(G4953GAT_1871_ngat) );
INVXL U_g4198 (.A(G4891GAT_1849_gat), .Y(G4891GAT_1849_ngat) );
INVXL U_g4199 (.A(G4950GAT_1873_gat), .Y(G4950GAT_1873_ngat) );
INVXL U_g4200 (.A(G4886GAT_1851_gat), .Y(G4886GAT_1851_ngat) );
INVXL U_g4201 (.A(G4947GAT_1875_gat), .Y(G4947GAT_1875_ngat) );
INVXL U_g4202 (.A(G4881GAT_1853_gat), .Y(G4881GAT_1853_ngat) );
INVXL U_g4203 (.A(G5063GAT_1879_gat), .Y(G5063GAT_1879_ngat) );
INVXL U_g4204 (.A(G5064GAT_1880_gat), .Y(G5064GAT_1880_ngat) );
INVXL U_g4205 (.A(G5059GAT_1881_gat), .Y(G5059GAT_1881_ngat) );
INVXL U_g4206 (.A(G5056GAT_1882_gat), .Y(G5056GAT_1882_ngat) );
INVXL U_g4207 (.A(G5053GAT_1883_gat), .Y(G5053GAT_1883_ngat) );
INVXL U_g4208 (.A(G5051GAT_1884_gat), .Y(G5051GAT_1884_ngat) );
INVXL U_g4209 (.A(G5052GAT_1894_gat), .Y(G5052GAT_1894_ngat) );
INVXL U_g4210 (.A(G5047GAT_1895_gat), .Y(G5047GAT_1895_ngat) );
INVXL U_g4211 (.A(G5042GAT_1886_gat), .Y(G5042GAT_1886_ngat) );
INVXL U_g4212 (.A(G5043GAT_1887_gat), .Y(G5043GAT_1887_ngat) );
INVXL U_g4213 (.A(G5038GAT_1888_gat), .Y(G5038GAT_1888_ngat) );
INVXL U_g4214 (.A(G5035GAT_1889_gat), .Y(G5035GAT_1889_ngat) );
INVXL U_g4215 (.A(G5032GAT_1890_gat), .Y(G5032GAT_1890_ngat) );
INVXL U_g4216 (.A(G5030GAT_1891_gat), .Y(G5030GAT_1891_ngat) );
INVXL U_g4217 (.A(G5031GAT_1896_gat), .Y(G5031GAT_1896_ngat) );
INVXL U_g4218 (.A(G5026GAT_1897_gat), .Y(G5026GAT_1897_ngat) );
INVXL U_g4219 (.A(G5021GAT_1893_gat), .Y(G5021GAT_1893_ngat) );
INVXL U_g4220 (.A(G5022GAT_1898_gat), .Y(G5022GAT_1898_ngat) );
INVXL U_g4221 (.A(G5017GAT_1899_gat), .Y(G5017GAT_1899_ngat) );
INVXL U_g4222 (.A(G5013GAT_1900_gat), .Y(G5013GAT_1900_ngat) );
INVXL U_g4223 (.A(G5009GAT_1901_gat), .Y(G5009GAT_1901_ngat) );
INVXL U_g4224 (.A(G5005GAT_1902_gat), .Y(G5005GAT_1902_ngat) );
INVXL U_g4225 (.A(G5044GAT_1885_gat), .Y(G5044GAT_1885_ngat) );
INVXL U_g4226 (.A(G1062GAT_114_gat), .Y(G1062GAT_114_ngat) );
INVXL U_g4227 (.A(G5023GAT_1892_gat), .Y(G5023GAT_1892_ngat) );
INVXL U_g4228 (.A(G819GAT_195_gat), .Y(G819GAT_195_ngat) );
INVXL U_g4229 (.A(G5113GAT_1904_gat), .Y(G5113GAT_1904_ngat) );
INVXL U_g4230 (.A(G5114GAT_1905_gat), .Y(G5114GAT_1905_ngat) );
INVXL U_g4231 (.A(G5109GAT_1906_gat), .Y(G5109GAT_1906_ngat) );
INVXL U_g4232 (.A(G5106GAT_1907_gat), .Y(G5106GAT_1907_ngat) );
INVXL U_g4233 (.A(G5103GAT_1908_gat), .Y(G5103GAT_1908_ngat) );
INVXL U_g4234 (.A(G5101GAT_1909_gat), .Y(G5101GAT_1909_ngat) );
INVXL U_g4235 (.A(G5102GAT_1922_gat), .Y(G5102GAT_1922_ngat) );
INVXL U_g4236 (.A(G5097GAT_1923_gat), .Y(G5097GAT_1923_ngat) );
INVXL U_g4237 (.A(G5092GAT_1911_gat), .Y(G5092GAT_1911_ngat) );
INVXL U_g4238 (.A(G5093GAT_1912_gat), .Y(G5093GAT_1912_ngat) );
INVXL U_g4239 (.A(G5088GAT_1913_gat), .Y(G5088GAT_1913_ngat) );
INVXL U_g4240 (.A(G5085GAT_1914_gat), .Y(G5085GAT_1914_ngat) );
INVXL U_g4241 (.A(G5082GAT_1915_gat), .Y(G5082GAT_1915_ngat) );
INVXL U_g4242 (.A(G5080GAT_1916_gat), .Y(G5080GAT_1916_ngat) );
INVXL U_g4243 (.A(G5081GAT_1924_gat), .Y(G5081GAT_1924_ngat) );
INVXL U_g4244 (.A(G5076GAT_1925_gat), .Y(G5076GAT_1925_ngat) );
INVXL U_g4245 (.A(G5071GAT_1918_gat), .Y(G5071GAT_1918_ngat) );
INVXL U_g4246 (.A(G5072GAT_1926_gat), .Y(G5072GAT_1926_ngat) );
INVXL U_g4247 (.A(G5115GAT_1903_gat), .Y(G5115GAT_1903_ngat) );
INVXL U_g4248 (.A(G1257GAT_49_gat), .Y(G1257GAT_49_ngat) );
INVXL U_g4249 (.A(G5069GAT_1919_gat), .Y(G5069GAT_1919_ngat) );
INVXL U_g4250 (.A(G5070GAT_1927_gat), .Y(G5070GAT_1927_ngat) );
INVXL U_g4251 (.A(G5067GAT_1920_gat), .Y(G5067GAT_1920_ngat) );
INVXL U_g4252 (.A(G5068GAT_1928_gat), .Y(G5068GAT_1928_ngat) );
INVXL U_g4253 (.A(G5065GAT_1921_gat), .Y(G5065GAT_1921_ngat) );
INVXL U_g4254 (.A(G5066GAT_1929_gat), .Y(G5066GAT_1929_ngat) );
INVXL U_g4255 (.A(G5094GAT_1910_gat), .Y(G5094GAT_1910_ngat) );
INVXL U_g4256 (.A(G1014GAT_130_gat), .Y(G1014GAT_130_ngat) );
INVXL U_g4257 (.A(G5073GAT_1917_gat), .Y(G5073GAT_1917_ngat) );
INVXL U_g4258 (.A(G771GAT_211_gat), .Y(G771GAT_211_ngat) );
INVXL U_g4259 (.A(G5172GAT_1945_gat), .Y(G5172GAT_1945_ngat) );
INVXL U_g4260 (.A(G5167GAT_1931_gat), .Y(G5167GAT_1931_ngat) );
INVXL U_g4261 (.A(G5168GAT_1932_gat), .Y(G5168GAT_1932_ngat) );
INVXL U_g4262 (.A(G5163GAT_1933_gat), .Y(G5163GAT_1933_ngat) );
INVXL U_g4263 (.A(G5160GAT_1934_gat), .Y(G5160GAT_1934_ngat) );
INVXL U_g4264 (.A(G5157GAT_1935_gat), .Y(G5157GAT_1935_ngat) );
INVXL U_g4265 (.A(G5155GAT_1936_gat), .Y(G5155GAT_1936_ngat) );
INVXL U_g4266 (.A(G5156GAT_1949_gat), .Y(G5156GAT_1949_ngat) );
INVXL U_g4267 (.A(G5151GAT_1950_gat), .Y(G5151GAT_1950_ngat) );
INVXL U_g4268 (.A(G5146GAT_1938_gat), .Y(G5146GAT_1938_ngat) );
INVXL U_g4269 (.A(G5147GAT_1939_gat), .Y(G5147GAT_1939_ngat) );
INVXL U_g4270 (.A(G5142GAT_1940_gat), .Y(G5142GAT_1940_ngat) );
INVXL U_g4271 (.A(G5139GAT_1941_gat), .Y(G5139GAT_1941_ngat) );
INVXL U_g4272 (.A(G5136GAT_1942_gat), .Y(G5136GAT_1942_ngat) );
INVXL U_g4273 (.A(G5134GAT_1943_gat), .Y(G5134GAT_1943_ngat) );
INVXL U_g4274 (.A(G5135GAT_1951_gat), .Y(G5135GAT_1951_ngat) );
INVXL U_g4275 (.A(G5130GAT_1952_gat), .Y(G5130GAT_1952_ngat) );
INVXL U_g4276 (.A(G5169GAT_1930_gat), .Y(G5169GAT_1930_ngat) );
INVXL U_g4277 (.A(G1209GAT_65_gat), .Y(G1209GAT_65_ngat) );
INVXL U_g4278 (.A(G5148GAT_1937_gat), .Y(G5148GAT_1937_ngat) );
INVXL U_g4279 (.A(G966GAT_146_gat), .Y(G966GAT_146_ngat) );
INVXL U_g4280 (.A(G5127GAT_1944_gat), .Y(G5127GAT_1944_ngat) );
INVXL U_g4281 (.A(G723GAT_227_gat), .Y(G723GAT_227_ngat) );
INVXL U_g4282 (.A(G5124GAT_1946_gat), .Y(G5124GAT_1946_ngat) );
INVXL U_g4283 (.A(G675GAT_243_gat), .Y(G675GAT_243_ngat) );
INVXL U_g4284 (.A(G5121GAT_1947_gat), .Y(G5121GAT_1947_ngat) );
INVXL U_g4285 (.A(G627GAT_259_gat), .Y(G627GAT_259_ngat) );
INVXL U_g4286 (.A(G5118GAT_1948_gat), .Y(G5118GAT_1948_ngat) );
INVXL U_g4287 (.A(G579GAT_275_gat), .Y(G579GAT_275_ngat) );
INVXL U_g4288 (.A(G1305GAT_33_gat), .Y(G1305GAT_33_ngat) );
INVXL U_g4289 (.A(G5236GAT_1953_gat), .Y(G5236GAT_1953_ngat) );
INVXL U_g4290 (.A(G5234GAT_1954_gat), .Y(G5234GAT_1954_ngat) );
INVXL U_g4291 (.A(G5235GAT_1969_gat), .Y(G5235GAT_1969_ngat) );
INVXL U_g4292 (.A(G5230GAT_1970_gat), .Y(G5230GAT_1970_ngat) );
INVXL U_g4293 (.A(G5225GAT_1956_gat), .Y(G5225GAT_1956_ngat) );
INVXL U_g4294 (.A(G5226GAT_1957_gat), .Y(G5226GAT_1957_ngat) );
INVXL U_g4295 (.A(G5221GAT_1958_gat), .Y(G5221GAT_1958_ngat) );
INVXL U_g4296 (.A(G5218GAT_1959_gat), .Y(G5218GAT_1959_ngat) );
INVXL U_g4297 (.A(G5215GAT_1960_gat), .Y(G5215GAT_1960_ngat) );
INVXL U_g4298 (.A(G5213GAT_1961_gat), .Y(G5213GAT_1961_ngat) );
INVXL U_g4299 (.A(G5214GAT_1971_gat), .Y(G5214GAT_1971_ngat) );
INVXL U_g4300 (.A(G5209GAT_1972_gat), .Y(G5209GAT_1972_ngat) );
INVXL U_g4301 (.A(G5204GAT_1963_gat), .Y(G5204GAT_1963_ngat) );
INVXL U_g4302 (.A(G5205GAT_1964_gat), .Y(G5205GAT_1964_ngat) );
INVXL U_g4303 (.A(G5200GAT_1965_gat), .Y(G5200GAT_1965_ngat) );
INVXL U_g4304 (.A(G5197GAT_1966_gat), .Y(G5197GAT_1966_ngat) );
INVXL U_g4305 (.A(G5194GAT_1967_gat), .Y(G5194GAT_1967_ngat) );
INVXL U_g4306 (.A(G5192GAT_1968_gat), .Y(G5192GAT_1968_ngat) );
INVXL U_g4307 (.A(G5193GAT_1973_gat), .Y(G5193GAT_1973_ngat) );
INVXL U_g4308 (.A(G5188GAT_1974_gat), .Y(G5188GAT_1974_ngat) );
INVXL U_g4309 (.A(G5184GAT_1975_gat), .Y(G5184GAT_1975_ngat) );
INVXL U_g4310 (.A(G5180GAT_1976_gat), .Y(G5180GAT_1976_ngat) );
INVXL U_g4311 (.A(G5227GAT_1955_gat), .Y(G5227GAT_1955_ngat) );
INVXL U_g4312 (.A(G1161GAT_81_gat), .Y(G1161GAT_81_ngat) );
INVXL U_g4313 (.A(G5176GAT_1977_gat), .Y(G5176GAT_1977_ngat) );
INVXL U_g4314 (.A(G5206GAT_1962_gat), .Y(G5206GAT_1962_ngat) );
INVXL U_g4315 (.A(G918GAT_162_gat), .Y(G918GAT_162_ngat) );
INVXL U_g4316 (.A(G5304GAT_1978_gat), .Y(G5304GAT_1978_ngat) );
INVXL U_g4317 (.A(G5301GAT_1979_gat), .Y(G5301GAT_1979_ngat) );
INVXL U_g4318 (.A(G5298GAT_1980_gat), .Y(G5298GAT_1980_ngat) );
INVXL U_g4319 (.A(G5296GAT_1981_gat), .Y(G5296GAT_1981_ngat) );
INVXL U_g4320 (.A(G5297GAT_1996_gat), .Y(G5297GAT_1996_ngat) );
INVXL U_g4321 (.A(G5292GAT_1998_gat), .Y(G5292GAT_1998_ngat) );
INVXL U_g4322 (.A(G5287GAT_1983_gat), .Y(G5287GAT_1983_ngat) );
INVXL U_g4323 (.A(G5288GAT_1984_gat), .Y(G5288GAT_1984_ngat) );
INVXL U_g4324 (.A(G5283GAT_1985_gat), .Y(G5283GAT_1985_ngat) );
INVXL U_g4325 (.A(G5280GAT_1986_gat), .Y(G5280GAT_1986_ngat) );
INVXL U_g4326 (.A(G5277GAT_1987_gat), .Y(G5277GAT_1987_ngat) );
INVXL U_g4327 (.A(G5275GAT_1988_gat), .Y(G5275GAT_1988_ngat) );
INVXL U_g4328 (.A(G5276GAT_2000_gat), .Y(G5276GAT_2000_ngat) );
INVXL U_g4329 (.A(G5271GAT_2001_gat), .Y(G5271GAT_2001_ngat) );
INVXL U_g4330 (.A(G5266GAT_1990_gat), .Y(G5266GAT_1990_ngat) );
INVXL U_g4331 (.A(G5267GAT_1991_gat), .Y(G5267GAT_1991_ngat) );
INVXL U_g4332 (.A(G5262GAT_1992_gat), .Y(G5262GAT_1992_ngat) );
INVXL U_g4333 (.A(G5259GAT_1993_gat), .Y(G5259GAT_1993_ngat) );
INVXL U_g4334 (.A(G5256GAT_2002_gat), .Y(G5256GAT_2002_ngat) );
INVXL U_g4335 (.A(G5254GAT_1994_gat), .Y(G5254GAT_1994_ngat) );
INVXL U_g4336 (.A(G5255GAT_2003_gat), .Y(G5255GAT_2003_ngat) );
INVXL U_g4337 (.A(G5249GAT_1995_gat), .Y(G5249GAT_1995_ngat) );
INVXL U_g4338 (.A(G5250GAT_2005_gat), .Y(G5250GAT_2005_ngat) );
INVXL U_g4339 (.A(G5244GAT_1997_gat), .Y(G5244GAT_1997_ngat) );
INVXL U_g4340 (.A(G5245GAT_2007_gat), .Y(G5245GAT_2007_ngat) );
INVXL U_g4341 (.A(G5239GAT_1999_gat), .Y(G5239GAT_1999_ngat) );
INVXL U_g4342 (.A(G5240GAT_2009_gat), .Y(G5240GAT_2009_ngat) );
INVXL U_g4343 (.A(G5289GAT_1982_gat), .Y(G5289GAT_1982_ngat) );
INVXL U_g4344 (.A(G1113GAT_97_gat), .Y(G1113GAT_97_ngat) );
INVXL U_g4345 (.A(G5268GAT_1989_gat), .Y(G5268GAT_1989_ngat) );
INVXL U_g4346 (.A(G870GAT_178_gat), .Y(G870GAT_178_ngat) );
INVXL U_g4347 (.A(G5364GAT_2010_gat), .Y(G5364GAT_2010_ngat) );
INVXL U_g4348 (.A(G5365GAT_2011_gat), .Y(G5365GAT_2011_ngat) );
INVXL U_g4349 (.A(G5360GAT_2012_gat), .Y(G5360GAT_2012_ngat) );
INVXL U_g4350 (.A(G5357GAT_2013_gat), .Y(G5357GAT_2013_ngat) );
INVXL U_g4351 (.A(G5354GAT_2014_gat), .Y(G5354GAT_2014_ngat) );
INVXL U_g4352 (.A(G5352GAT_2015_gat), .Y(G5352GAT_2015_ngat) );
INVXL U_g4353 (.A(G5353GAT_2030_gat), .Y(G5353GAT_2030_ngat) );
INVXL U_g4354 (.A(G5348GAT_2032_gat), .Y(G5348GAT_2032_ngat) );
INVXL U_g4355 (.A(G5343GAT_2017_gat), .Y(G5343GAT_2017_ngat) );
INVXL U_g4356 (.A(G5344GAT_2018_gat), .Y(G5344GAT_2018_ngat) );
INVXL U_g4357 (.A(G5339GAT_2019_gat), .Y(G5339GAT_2019_ngat) );
INVXL U_g4358 (.A(G5336GAT_2020_gat), .Y(G5336GAT_2020_ngat) );
INVXL U_g4359 (.A(G5333GAT_2021_gat), .Y(G5333GAT_2021_ngat) );
INVXL U_g4360 (.A(G5331GAT_2022_gat), .Y(G5331GAT_2022_ngat) );
INVXL U_g4361 (.A(G5332GAT_2033_gat), .Y(G5332GAT_2033_ngat) );
INVXL U_g4362 (.A(G5327GAT_2034_gat), .Y(G5327GAT_2034_ngat) );
INVXL U_g4363 (.A(G5322GAT_2024_gat), .Y(G5322GAT_2024_ngat) );
INVXL U_g4364 (.A(G5323GAT_2025_gat), .Y(G5323GAT_2025_ngat) );
INVXL U_g4365 (.A(G5318GAT_2026_gat), .Y(G5318GAT_2026_ngat) );
INVXL U_g4366 (.A(G5345GAT_2016_gat), .Y(G5345GAT_2016_ngat) );
INVXL U_g4367 (.A(G1065GAT_113_gat), .Y(G1065GAT_113_ngat) );
INVXL U_g4368 (.A(G5324GAT_2023_gat), .Y(G5324GAT_2023_ngat) );
INVXL U_g4369 (.A(G822GAT_194_gat), .Y(G822GAT_194_ngat) );
INVXL U_g4370 (.A(G5315GAT_2027_gat), .Y(G5315GAT_2027_ngat) );
INVXL U_g4371 (.A(G5251GAT_2004_gat), .Y(G5251GAT_2004_ngat) );
INVXL U_g4372 (.A(G5312GAT_2028_gat), .Y(G5312GAT_2028_ngat) );
INVXL U_g4373 (.A(G5246GAT_2006_gat), .Y(G5246GAT_2006_ngat) );
INVXL U_g4374 (.A(G5309GAT_2029_gat), .Y(G5309GAT_2029_ngat) );
INVXL U_g4375 (.A(G5241GAT_2008_gat), .Y(G5241GAT_2008_ngat) );
INVXL U_g4376 (.A(G5420GAT_2036_gat), .Y(G5420GAT_2036_ngat) );
INVXL U_g4377 (.A(G5421GAT_2037_gat), .Y(G5421GAT_2037_ngat) );
INVXL U_g4378 (.A(G5416GAT_2038_gat), .Y(G5416GAT_2038_ngat) );
INVXL U_g4379 (.A(G5413GAT_2039_gat), .Y(G5413GAT_2039_ngat) );
INVXL U_g4380 (.A(G5410GAT_2040_gat), .Y(G5410GAT_2040_ngat) );
INVXL U_g4381 (.A(G5408GAT_2041_gat), .Y(G5408GAT_2041_ngat) );
INVXL U_g4382 (.A(G5409GAT_2051_gat), .Y(G5409GAT_2051_ngat) );
INVXL U_g4383 (.A(G5404GAT_2052_gat), .Y(G5404GAT_2052_ngat) );
INVXL U_g4384 (.A(G5399GAT_2043_gat), .Y(G5399GAT_2043_ngat) );
INVXL U_g4385 (.A(G5400GAT_2044_gat), .Y(G5400GAT_2044_ngat) );
INVXL U_g4386 (.A(G5395GAT_2045_gat), .Y(G5395GAT_2045_ngat) );
INVXL U_g4387 (.A(G5392GAT_2046_gat), .Y(G5392GAT_2046_ngat) );
INVXL U_g4388 (.A(G5389GAT_2047_gat), .Y(G5389GAT_2047_ngat) );
INVXL U_g4389 (.A(G5387GAT_2048_gat), .Y(G5387GAT_2048_ngat) );
INVXL U_g4390 (.A(G5388GAT_2053_gat), .Y(G5388GAT_2053_ngat) );
INVXL U_g4391 (.A(G5383GAT_2054_gat), .Y(G5383GAT_2054_ngat) );
INVXL U_g4392 (.A(G5378GAT_2050_gat), .Y(G5378GAT_2050_ngat) );
INVXL U_g4393 (.A(G5379GAT_2055_gat), .Y(G5379GAT_2055_ngat) );
INVXL U_g4394 (.A(G5374GAT_2056_gat), .Y(G5374GAT_2056_ngat) );
INVXL U_g4395 (.A(G5422GAT_2035_gat), .Y(G5422GAT_2035_ngat) );
INVXL U_g4396 (.A(G1260GAT_48_gat), .Y(G1260GAT_48_ngat) );
INVXL U_g4397 (.A(G5370GAT_2057_gat), .Y(G5370GAT_2057_ngat) );
INVXL U_g4398 (.A(G5366GAT_2058_gat), .Y(G5366GAT_2058_ngat) );
INVXL U_g4399 (.A(G5401GAT_2042_gat), .Y(G5401GAT_2042_ngat) );
INVXL U_g4400 (.A(G1017GAT_129_gat), .Y(G1017GAT_129_ngat) );
INVXL U_g4401 (.A(G5380GAT_2049_gat), .Y(G5380GAT_2049_ngat) );
INVXL U_g4402 (.A(G774GAT_210_gat), .Y(G774GAT_210_ngat) );
INVXL U_g4403 (.A(G5476GAT_2075_gat), .Y(G5476GAT_2075_ngat) );
INVXL U_g4404 (.A(G5471GAT_2060_gat), .Y(G5471GAT_2060_ngat) );
INVXL U_g4405 (.A(G5472GAT_2061_gat), .Y(G5472GAT_2061_ngat) );
INVXL U_g4406 (.A(G5467GAT_2062_gat), .Y(G5467GAT_2062_ngat) );
INVXL U_g4407 (.A(G5464GAT_2063_gat), .Y(G5464GAT_2063_ngat) );
INVXL U_g4408 (.A(G5461GAT_2064_gat), .Y(G5461GAT_2064_ngat) );
INVXL U_g4409 (.A(G5459GAT_2065_gat), .Y(G5459GAT_2065_ngat) );
INVXL U_g4410 (.A(G5460GAT_2078_gat), .Y(G5460GAT_2078_ngat) );
INVXL U_g4411 (.A(G5455GAT_2079_gat), .Y(G5455GAT_2079_ngat) );
INVXL U_g4412 (.A(G5450GAT_2067_gat), .Y(G5450GAT_2067_ngat) );
INVXL U_g4413 (.A(G5451GAT_2068_gat), .Y(G5451GAT_2068_ngat) );
INVXL U_g4414 (.A(G5446GAT_2069_gat), .Y(G5446GAT_2069_ngat) );
INVXL U_g4415 (.A(G5443GAT_2070_gat), .Y(G5443GAT_2070_ngat) );
INVXL U_g4416 (.A(G5440GAT_2071_gat), .Y(G5440GAT_2071_ngat) );
INVXL U_g4417 (.A(G5438GAT_2072_gat), .Y(G5438GAT_2072_ngat) );
INVXL U_g4418 (.A(G5439GAT_2080_gat), .Y(G5439GAT_2080_ngat) );
INVXL U_g4419 (.A(G5434GAT_2081_gat), .Y(G5434GAT_2081_ngat) );
INVXL U_g4420 (.A(G5429GAT_2074_gat), .Y(G5429GAT_2074_ngat) );
INVXL U_g4421 (.A(G5430GAT_2082_gat), .Y(G5430GAT_2082_ngat) );
INVXL U_g4422 (.A(G5427GAT_2076_gat), .Y(G5427GAT_2076_ngat) );
INVXL U_g4423 (.A(G5428GAT_2083_gat), .Y(G5428GAT_2083_ngat) );
INVXL U_g4424 (.A(G5473GAT_2059_gat), .Y(G5473GAT_2059_ngat) );
INVXL U_g4425 (.A(G1212GAT_64_gat), .Y(G1212GAT_64_ngat) );
INVXL U_g4426 (.A(G5425GAT_2077_gat), .Y(G5425GAT_2077_ngat) );
INVXL U_g4427 (.A(G5426GAT_2084_gat), .Y(G5426GAT_2084_ngat) );
INVXL U_g4428 (.A(G5452GAT_2066_gat), .Y(G5452GAT_2066_ngat) );
INVXL U_g4429 (.A(G969GAT_145_gat), .Y(G969GAT_145_ngat) );
INVXL U_g4430 (.A(G5431GAT_2073_gat), .Y(G5431GAT_2073_ngat) );
INVXL U_g4431 (.A(G726GAT_226_gat), .Y(G726GAT_226_ngat) );
INVXL U_g4432 (.A(G1308GAT_32_gat), .Y(G1308GAT_32_ngat) );
INVXL U_g4433 (.A(G5537GAT_2085_gat), .Y(G5537GAT_2085_ngat) );
INVXL U_g4434 (.A(G5535GAT_2086_gat), .Y(G5535GAT_2086_ngat) );
INVXL U_g4435 (.A(G5536GAT_2102_gat), .Y(G5536GAT_2102_ngat) );
INVXL U_g4436 (.A(G5531GAT_2104_gat), .Y(G5531GAT_2104_ngat) );
INVXL U_g4437 (.A(G5526GAT_2088_gat), .Y(G5526GAT_2088_ngat) );
INVXL U_g4438 (.A(G5527GAT_2089_gat), .Y(G5527GAT_2089_ngat) );
INVXL U_g4439 (.A(G5522GAT_2090_gat), .Y(G5522GAT_2090_ngat) );
INVXL U_g4440 (.A(G5519GAT_2091_gat), .Y(G5519GAT_2091_ngat) );
INVXL U_g4441 (.A(G5516GAT_2092_gat), .Y(G5516GAT_2092_ngat) );
INVXL U_g4442 (.A(G5514GAT_2093_gat), .Y(G5514GAT_2093_ngat) );
INVXL U_g4443 (.A(G5515GAT_2106_gat), .Y(G5515GAT_2106_ngat) );
INVXL U_g4444 (.A(G5510GAT_2107_gat), .Y(G5510GAT_2107_ngat) );
INVXL U_g4445 (.A(G5505GAT_2095_gat), .Y(G5505GAT_2095_ngat) );
INVXL U_g4446 (.A(G5506GAT_2096_gat), .Y(G5506GAT_2096_ngat) );
INVXL U_g4447 (.A(G5501GAT_2097_gat), .Y(G5501GAT_2097_ngat) );
INVXL U_g4448 (.A(G5498GAT_2098_gat), .Y(G5498GAT_2098_ngat) );
INVXL U_g4449 (.A(G5495GAT_2099_gat), .Y(G5495GAT_2099_ngat) );
INVXL U_g4450 (.A(G5493GAT_2100_gat), .Y(G5493GAT_2100_ngat) );
INVXL U_g4451 (.A(G5494GAT_2108_gat), .Y(G5494GAT_2108_ngat) );
INVXL U_g4452 (.A(G5489GAT_2109_gat), .Y(G5489GAT_2109_ngat) );
INVXL U_g4453 (.A(G5528GAT_2087_gat), .Y(G5528GAT_2087_ngat) );
INVXL U_g4454 (.A(G1164GAT_80_gat), .Y(G1164GAT_80_ngat) );
INVXL U_g4455 (.A(G5507GAT_2094_gat), .Y(G5507GAT_2094_ngat) );
INVXL U_g4456 (.A(G921GAT_161_gat), .Y(G921GAT_161_ngat) );
INVXL U_g4457 (.A(G5486GAT_2101_gat), .Y(G5486GAT_2101_ngat) );
INVXL U_g4458 (.A(G678GAT_242_gat), .Y(G678GAT_242_ngat) );
INVXL U_g4459 (.A(G5483GAT_2103_gat), .Y(G5483GAT_2103_ngat) );
INVXL U_g4460 (.A(G630GAT_258_gat), .Y(G630GAT_258_ngat) );
INVXL U_g4461 (.A(G5480GAT_2105_gat), .Y(G5480GAT_2105_ngat) );
INVXL U_g4462 (.A(G582GAT_274_gat), .Y(G582GAT_274_ngat) );
INVXL U_g4463 (.A(G5602GAT_2110_gat), .Y(G5602GAT_2110_ngat) );
INVXL U_g4464 (.A(G5599GAT_2111_gat), .Y(G5599GAT_2111_ngat) );
INVXL U_g4465 (.A(G5596GAT_2112_gat), .Y(G5596GAT_2112_ngat) );
INVXL U_g4466 (.A(G5594GAT_2113_gat), .Y(G5594GAT_2113_ngat) );
INVXL U_g4467 (.A(G5595GAT_2128_gat), .Y(G5595GAT_2128_ngat) );
INVXL U_g4468 (.A(G5590GAT_2129_gat), .Y(G5590GAT_2129_ngat) );
INVXL U_g4469 (.A(G5585GAT_2115_gat), .Y(G5585GAT_2115_ngat) );
INVXL U_g4470 (.A(G5586GAT_2116_gat), .Y(G5586GAT_2116_ngat) );
INVXL U_g4471 (.A(G5581GAT_2117_gat), .Y(G5581GAT_2117_ngat) );
INVXL U_g4472 (.A(G5578GAT_2118_gat), .Y(G5578GAT_2118_ngat) );
INVXL U_g4473 (.A(G5575GAT_2119_gat), .Y(G5575GAT_2119_ngat) );
INVXL U_g4474 (.A(G5573GAT_2120_gat), .Y(G5573GAT_2120_ngat) );
INVXL U_g4475 (.A(G5574GAT_2130_gat), .Y(G5574GAT_2130_ngat) );
INVXL U_g4476 (.A(G5569GAT_2131_gat), .Y(G5569GAT_2131_ngat) );
INVXL U_g4477 (.A(G5564GAT_2122_gat), .Y(G5564GAT_2122_ngat) );
INVXL U_g4478 (.A(G5565GAT_2123_gat), .Y(G5565GAT_2123_ngat) );
INVXL U_g4479 (.A(G5560GAT_2124_gat), .Y(G5560GAT_2124_ngat) );
INVXL U_g4480 (.A(G5557GAT_2125_gat), .Y(G5557GAT_2125_ngat) );
INVXL U_g4481 (.A(G5554GAT_2126_gat), .Y(G5554GAT_2126_ngat) );
INVXL U_g4482 (.A(G5552GAT_2127_gat), .Y(G5552GAT_2127_ngat) );
INVXL U_g4483 (.A(G5553GAT_2132_gat), .Y(G5553GAT_2132_ngat) );
INVXL U_g4484 (.A(G5548GAT_2133_gat), .Y(G5548GAT_2133_ngat) );
INVXL U_g4485 (.A(G5544GAT_2134_gat), .Y(G5544GAT_2134_ngat) );
INVXL U_g4486 (.A(G5540GAT_2135_gat), .Y(G5540GAT_2135_ngat) );
INVXL U_g4487 (.A(G5587GAT_2114_gat), .Y(G5587GAT_2114_ngat) );
INVXL U_g4488 (.A(G1116GAT_96_gat), .Y(G1116GAT_96_ngat) );
INVXL U_g4489 (.A(G5566GAT_2121_gat), .Y(G5566GAT_2121_ngat) );
INVXL U_g4490 (.A(G873GAT_177_gat), .Y(G873GAT_177_ngat) );
INVXL U_g4491 (.A(G5670GAT_2136_gat), .Y(G5670GAT_2136_ngat) );
INVXL U_g4492 (.A(G5671GAT_2137_gat), .Y(G5671GAT_2137_ngat) );
INVXL U_g4493 (.A(G5666GAT_2138_gat), .Y(G5666GAT_2138_ngat) );
INVXL U_g4494 (.A(G5663GAT_2139_gat), .Y(G5663GAT_2139_ngat) );
INVXL U_g4495 (.A(G5660GAT_2140_gat), .Y(G5660GAT_2140_ngat) );
INVXL U_g4496 (.A(G5658GAT_2141_gat), .Y(G5658GAT_2141_ngat) );
INVXL U_g4497 (.A(G5659GAT_2157_gat), .Y(G5659GAT_2157_ngat) );
INVXL U_g4498 (.A(G5654GAT_2158_gat), .Y(G5654GAT_2158_ngat) );
INVXL U_g4499 (.A(G5649GAT_2143_gat), .Y(G5649GAT_2143_ngat) );
INVXL U_g4500 (.A(G5650GAT_2144_gat), .Y(G5650GAT_2144_ngat) );
INVXL U_g4501 (.A(G5645GAT_2145_gat), .Y(G5645GAT_2145_ngat) );
INVXL U_g4502 (.A(G5642GAT_2146_gat), .Y(G5642GAT_2146_ngat) );
INVXL U_g4503 (.A(G5639GAT_2147_gat), .Y(G5639GAT_2147_ngat) );
INVXL U_g4504 (.A(G5637GAT_2148_gat), .Y(G5637GAT_2148_ngat) );
INVXL U_g4505 (.A(G5638GAT_2159_gat), .Y(G5638GAT_2159_ngat) );
INVXL U_g4506 (.A(G5633GAT_2160_gat), .Y(G5633GAT_2160_ngat) );
INVXL U_g4507 (.A(G5628GAT_2150_gat), .Y(G5628GAT_2150_ngat) );
INVXL U_g4508 (.A(G5629GAT_2151_gat), .Y(G5629GAT_2151_ngat) );
INVXL U_g4509 (.A(G5624GAT_2152_gat), .Y(G5624GAT_2152_ngat) );
INVXL U_g4510 (.A(G5621GAT_2153_gat), .Y(G5621GAT_2153_ngat) );
INVXL U_g4511 (.A(G5618GAT_2161_gat), .Y(G5618GAT_2161_ngat) );
INVXL U_g4512 (.A(G5616GAT_2154_gat), .Y(G5616GAT_2154_ngat) );
INVXL U_g4513 (.A(G5617GAT_2162_gat), .Y(G5617GAT_2162_ngat) );
INVXL U_g4514 (.A(G5611GAT_2155_gat), .Y(G5611GAT_2155_ngat) );
INVXL U_g4515 (.A(G5612GAT_2164_gat), .Y(G5612GAT_2164_ngat) );
INVXL U_g4516 (.A(G5606GAT_2156_gat), .Y(G5606GAT_2156_ngat) );
INVXL U_g4517 (.A(G5607GAT_2166_gat), .Y(G5607GAT_2166_ngat) );
INVXL U_g4518 (.A(G5651GAT_2142_gat), .Y(G5651GAT_2142_ngat) );
INVXL U_g4519 (.A(G1068GAT_112_gat), .Y(G1068GAT_112_ngat) );
INVXL U_g4520 (.A(G5630GAT_2149_gat), .Y(G5630GAT_2149_ngat) );
INVXL U_g4521 (.A(G825GAT_193_gat), .Y(G825GAT_193_ngat) );
INVXL U_g4522 (.A(G5725GAT_2168_gat), .Y(G5725GAT_2168_ngat) );
INVXL U_g4523 (.A(G5726GAT_2169_gat), .Y(G5726GAT_2169_ngat) );
INVXL U_g4524 (.A(G5721GAT_2170_gat), .Y(G5721GAT_2170_ngat) );
INVXL U_g4525 (.A(G5718GAT_2171_gat), .Y(G5718GAT_2171_ngat) );
INVXL U_g4526 (.A(G5715GAT_2172_gat), .Y(G5715GAT_2172_ngat) );
INVXL U_g4527 (.A(G5713GAT_2173_gat), .Y(G5713GAT_2173_ngat) );
INVXL U_g4528 (.A(G5714GAT_2188_gat), .Y(G5714GAT_2188_ngat) );
INVXL U_g4529 (.A(G5709GAT_2189_gat), .Y(G5709GAT_2189_ngat) );
INVXL U_g4530 (.A(G5704GAT_2175_gat), .Y(G5704GAT_2175_ngat) );
INVXL U_g4531 (.A(G5705GAT_2176_gat), .Y(G5705GAT_2176_ngat) );
INVXL U_g4532 (.A(G5700GAT_2177_gat), .Y(G5700GAT_2177_ngat) );
INVXL U_g4533 (.A(G5697GAT_2178_gat), .Y(G5697GAT_2178_ngat) );
INVXL U_g4534 (.A(G5694GAT_2179_gat), .Y(G5694GAT_2179_ngat) );
INVXL U_g4535 (.A(G5692GAT_2180_gat), .Y(G5692GAT_2180_ngat) );
INVXL U_g4536 (.A(G5693GAT_2190_gat), .Y(G5693GAT_2190_ngat) );
INVXL U_g4537 (.A(G5688GAT_2191_gat), .Y(G5688GAT_2191_ngat) );
INVXL U_g4538 (.A(G5683GAT_2182_gat), .Y(G5683GAT_2182_ngat) );
INVXL U_g4539 (.A(G5684GAT_2183_gat), .Y(G5684GAT_2183_ngat) );
INVXL U_g4540 (.A(G5679GAT_2184_gat), .Y(G5679GAT_2184_ngat) );
INVXL U_g4541 (.A(G5706GAT_2174_gat), .Y(G5706GAT_2174_ngat) );
INVXL U_g4542 (.A(G1020GAT_128_gat), .Y(G1020GAT_128_ngat) );
INVXL U_g4543 (.A(G5685GAT_2181_gat), .Y(G5685GAT_2181_ngat) );
INVXL U_g4544 (.A(G777GAT_209_gat), .Y(G777GAT_209_ngat) );
INVXL U_g4545 (.A(G5676GAT_2185_gat), .Y(G5676GAT_2185_ngat) );
INVXL U_g4546 (.A(G5613GAT_2163_gat), .Y(G5613GAT_2163_ngat) );
INVXL U_g4547 (.A(G5673GAT_2186_gat), .Y(G5673GAT_2186_ngat) );
INVXL U_g4548 (.A(G5608GAT_2165_gat), .Y(G5608GAT_2165_ngat) );
INVXL U_g4549 (.A(G5780GAT_2193_gat), .Y(G5780GAT_2193_ngat) );
INVXL U_g4550 (.A(G5781GAT_2194_gat), .Y(G5781GAT_2194_ngat) );
INVXL U_g4551 (.A(G5776GAT_2195_gat), .Y(G5776GAT_2195_ngat) );
INVXL U_g4552 (.A(G5773GAT_2196_gat), .Y(G5773GAT_2196_ngat) );
INVXL U_g4553 (.A(G5770GAT_2197_gat), .Y(G5770GAT_2197_ngat) );
INVXL U_g4554 (.A(G5768GAT_2198_gat), .Y(G5768GAT_2198_ngat) );
INVXL U_g4555 (.A(G5769GAT_2208_gat), .Y(G5769GAT_2208_ngat) );
INVXL U_g4556 (.A(G5764GAT_2209_gat), .Y(G5764GAT_2209_ngat) );
INVXL U_g4557 (.A(G5759GAT_2200_gat), .Y(G5759GAT_2200_ngat) );
INVXL U_g4558 (.A(G5760GAT_2201_gat), .Y(G5760GAT_2201_ngat) );
INVXL U_g4559 (.A(G5755GAT_2202_gat), .Y(G5755GAT_2202_ngat) );
INVXL U_g4560 (.A(G5752GAT_2203_gat), .Y(G5752GAT_2203_ngat) );
INVXL U_g4561 (.A(G5749GAT_2204_gat), .Y(G5749GAT_2204_ngat) );
INVXL U_g4562 (.A(G5747GAT_2205_gat), .Y(G5747GAT_2205_ngat) );
INVXL U_g4563 (.A(G5748GAT_2210_gat), .Y(G5748GAT_2210_ngat) );
INVXL U_g4564 (.A(G5743GAT_2211_gat), .Y(G5743GAT_2211_ngat) );
INVXL U_g4565 (.A(G5738GAT_2207_gat), .Y(G5738GAT_2207_ngat) );
INVXL U_g4566 (.A(G5739GAT_2212_gat), .Y(G5739GAT_2212_ngat) );
INVXL U_g4567 (.A(G5734GAT_2213_gat), .Y(G5734GAT_2213_ngat) );
INVXL U_g4568 (.A(G5730GAT_2214_gat), .Y(G5730GAT_2214_ngat) );
INVXL U_g4569 (.A(G5761GAT_2199_gat), .Y(G5761GAT_2199_ngat) );
INVXL U_g4570 (.A(G972GAT_144_gat), .Y(G972GAT_144_ngat) );
INVXL U_g4571 (.A(G5740GAT_2206_gat), .Y(G5740GAT_2206_ngat) );
INVXL U_g4572 (.A(G729GAT_225_gat), .Y(G729GAT_225_ngat) );
INVXL U_g4573 (.A(G5829GAT_2216_gat), .Y(G5829GAT_2216_ngat) );
INVXL U_g4574 (.A(G5830GAT_2217_gat), .Y(G5830GAT_2217_ngat) );
INVXL U_g4575 (.A(G5825GAT_2218_gat), .Y(G5825GAT_2218_ngat) );
INVXL U_g4576 (.A(G5822GAT_2219_gat), .Y(G5822GAT_2219_ngat) );
INVXL U_g4577 (.A(G5819GAT_2220_gat), .Y(G5819GAT_2220_ngat) );
INVXL U_g4578 (.A(G5817GAT_2221_gat), .Y(G5817GAT_2221_ngat) );
INVXL U_g4579 (.A(G5818GAT_2232_gat), .Y(G5818GAT_2232_ngat) );
INVXL U_g4580 (.A(G5813GAT_2233_gat), .Y(G5813GAT_2233_ngat) );
INVXL U_g4581 (.A(G5808GAT_2223_gat), .Y(G5808GAT_2223_ngat) );
INVXL U_g4582 (.A(G5809GAT_2224_gat), .Y(G5809GAT_2224_ngat) );
INVXL U_g4583 (.A(G5804GAT_2225_gat), .Y(G5804GAT_2225_ngat) );
INVXL U_g4584 (.A(G5801GAT_2226_gat), .Y(G5801GAT_2226_ngat) );
INVXL U_g4585 (.A(G5798GAT_2227_gat), .Y(G5798GAT_2227_ngat) );
INVXL U_g4586 (.A(G5796GAT_2228_gat), .Y(G5796GAT_2228_ngat) );
INVXL U_g4587 (.A(G5797GAT_2234_gat), .Y(G5797GAT_2234_ngat) );
INVXL U_g4588 (.A(G5792GAT_2235_gat), .Y(G5792GAT_2235_ngat) );
INVXL U_g4589 (.A(G5787GAT_2230_gat), .Y(G5787GAT_2230_ngat) );
INVXL U_g4590 (.A(G5788GAT_2236_gat), .Y(G5788GAT_2236_ngat) );
INVXL U_g4591 (.A(G5785GAT_2231_gat), .Y(G5785GAT_2231_ngat) );
INVXL U_g4592 (.A(G5786GAT_2237_gat), .Y(G5786GAT_2237_ngat) );
INVXL U_g4593 (.A(G5810GAT_2222_gat), .Y(G5810GAT_2222_ngat) );
INVXL U_g4594 (.A(G924GAT_160_gat), .Y(G924GAT_160_ngat) );
INVXL U_g4595 (.A(G5789GAT_2229_gat), .Y(G5789GAT_2229_ngat) );
INVXL U_g4596 (.A(G681GAT_241_gat), .Y(G681GAT_241_ngat) );
INVXL U_g4597 (.A(G5877GAT_2239_gat), .Y(G5877GAT_2239_ngat) );
INVXL U_g4598 (.A(G5878GAT_2240_gat), .Y(G5878GAT_2240_ngat) );
INVXL U_g4599 (.A(G5873GAT_2241_gat), .Y(G5873GAT_2241_ngat) );
INVXL U_g4600 (.A(G5870GAT_2242_gat), .Y(G5870GAT_2242_ngat) );
INVXL U_g4601 (.A(G5867GAT_2243_gat), .Y(G5867GAT_2243_ngat) );
INVXL U_g4602 (.A(G5865GAT_2244_gat), .Y(G5865GAT_2244_ngat) );
INVXL U_g4603 (.A(G5866GAT_2254_gat), .Y(G5866GAT_2254_ngat) );
INVXL U_g4604 (.A(G5861GAT_2255_gat), .Y(G5861GAT_2255_ngat) );
INVXL U_g4605 (.A(G5856GAT_2246_gat), .Y(G5856GAT_2246_ngat) );
INVXL U_g4606 (.A(G5857GAT_2247_gat), .Y(G5857GAT_2247_ngat) );
INVXL U_g4607 (.A(G5852GAT_2248_gat), .Y(G5852GAT_2248_ngat) );
INVXL U_g4608 (.A(G5849GAT_2249_gat), .Y(G5849GAT_2249_ngat) );
INVXL U_g4609 (.A(G5846GAT_2250_gat), .Y(G5846GAT_2250_ngat) );
INVXL U_g4610 (.A(G5844GAT_2251_gat), .Y(G5844GAT_2251_ngat) );
INVXL U_g4611 (.A(G5845GAT_2256_gat), .Y(G5845GAT_2256_ngat) );
INVXL U_g4612 (.A(G5840GAT_2257_gat), .Y(G5840GAT_2257_ngat) );
INVXL U_g4613 (.A(G5858GAT_2245_gat), .Y(G5858GAT_2245_ngat) );
INVXL U_g4614 (.A(G876GAT_176_gat), .Y(G876GAT_176_ngat) );
INVXL U_g4615 (.A(G5837GAT_2252_gat), .Y(G5837GAT_2252_ngat) );
INVXL U_g4616 (.A(G633GAT_257_gat), .Y(G633GAT_257_ngat) );
INVXL U_g4617 (.A(G5834GAT_2253_gat), .Y(G5834GAT_2253_ngat) );
INVXL U_g4618 (.A(G585GAT_273_gat), .Y(G585GAT_273_ngat) );
INVXL U_g4619 (.A(G5923GAT_2259_gat), .Y(G5923GAT_2259_ngat) );
INVXL U_g4620 (.A(G5924GAT_2260_gat), .Y(G5924GAT_2260_ngat) );
INVXL U_g4621 (.A(G5919GAT_2261_gat), .Y(G5919GAT_2261_ngat) );
INVXL U_g4622 (.A(G5916GAT_2262_gat), .Y(G5916GAT_2262_ngat) );
INVXL U_g4623 (.A(G5913GAT_2263_gat), .Y(G5913GAT_2263_ngat) );
INVXL U_g4624 (.A(G5911GAT_2264_gat), .Y(G5911GAT_2264_ngat) );
INVXL U_g4625 (.A(G5912GAT_2272_gat), .Y(G5912GAT_2272_ngat) );
INVXL U_g4626 (.A(G5907GAT_2273_gat), .Y(G5907GAT_2273_ngat) );
INVXL U_g4627 (.A(G5902GAT_2266_gat), .Y(G5902GAT_2266_ngat) );
INVXL U_g4628 (.A(G5903GAT_2267_gat), .Y(G5903GAT_2267_ngat) );
INVXL U_g4629 (.A(G5898GAT_2268_gat), .Y(G5898GAT_2268_ngat) );
INVXL U_g4630 (.A(G5895GAT_2269_gat), .Y(G5895GAT_2269_ngat) );
INVXL U_g4631 (.A(G5892GAT_2270_gat), .Y(G5892GAT_2270_ngat) );
INVXL U_g4632 (.A(G5890GAT_2271_gat), .Y(G5890GAT_2271_ngat) );
INVXL U_g4633 (.A(G5891GAT_2274_gat), .Y(G5891GAT_2274_ngat) );
INVXL U_g4634 (.A(G5886GAT_2275_gat), .Y(G5886GAT_2275_ngat) );
INVXL U_g4635 (.A(G5882GAT_2276_gat), .Y(G5882GAT_2276_ngat) );
INVXL U_g4636 (.A(G5904GAT_2265_gat), .Y(G5904GAT_2265_ngat) );
INVXL U_g4637 (.A(G828GAT_192_gat), .Y(G828GAT_192_ngat) );
INVXL U_g4638 (.A(G5966GAT_2278_gat), .Y(G5966GAT_2278_ngat) );
INVXL U_g4639 (.A(G5967GAT_2279_gat), .Y(G5967GAT_2279_ngat) );
INVXL U_g4640 (.A(G5962GAT_2280_gat), .Y(G5962GAT_2280_ngat) );
INVXL U_g4641 (.A(G5959GAT_2281_gat), .Y(G5959GAT_2281_ngat) );
INVXL U_g4642 (.A(G5956GAT_2282_gat), .Y(G5956GAT_2282_ngat) );
INVXL U_g4643 (.A(G5954GAT_2283_gat), .Y(G5954GAT_2283_ngat) );
INVXL U_g4644 (.A(G5955GAT_2291_gat), .Y(G5955GAT_2291_ngat) );
INVXL U_g4645 (.A(G5950GAT_2292_gat), .Y(G5950GAT_2292_ngat) );
INVXL U_g4646 (.A(G5945GAT_2285_gat), .Y(G5945GAT_2285_ngat) );
INVXL U_g4647 (.A(G5946GAT_2286_gat), .Y(G5946GAT_2286_ngat) );
INVXL U_g4648 (.A(G5941GAT_2287_gat), .Y(G5941GAT_2287_ngat) );
INVXL U_g4649 (.A(G5938GAT_2288_gat), .Y(G5938GAT_2288_ngat) );
INVXL U_g4650 (.A(G5935GAT_2293_gat), .Y(G5935GAT_2293_ngat) );
INVXL U_g4651 (.A(G5933GAT_2289_gat), .Y(G5933GAT_2289_ngat) );
INVXL U_g4652 (.A(G5934GAT_2294_gat), .Y(G5934GAT_2294_ngat) );
INVXL U_g4653 (.A(G5928GAT_2290_gat), .Y(G5928GAT_2290_ngat) );
INVXL U_g4654 (.A(G5929GAT_2296_gat), .Y(G5929GAT_2296_ngat) );
INVXL U_g4655 (.A(G5947GAT_2284_gat), .Y(G5947GAT_2284_ngat) );
INVXL U_g4656 (.A(G780GAT_208_gat), .Y(G780GAT_208_ngat) );
INVXL U_g4657 (.A(G6000GAT_2298_gat), .Y(G6000GAT_2298_ngat) );
INVXL U_g4658 (.A(G6001GAT_2299_gat), .Y(G6001GAT_2299_ngat) );
INVXL U_g4659 (.A(G5996GAT_2300_gat), .Y(G5996GAT_2300_ngat) );
INVXL U_g4660 (.A(G5993GAT_2301_gat), .Y(G5993GAT_2301_ngat) );
INVXL U_g4661 (.A(G5990GAT_2302_gat), .Y(G5990GAT_2302_ngat) );
INVXL U_g4662 (.A(G5988GAT_2303_gat), .Y(G5988GAT_2303_ngat) );
INVXL U_g4663 (.A(G5989GAT_2310_gat), .Y(G5989GAT_2310_ngat) );
INVXL U_g4664 (.A(G5984GAT_2311_gat), .Y(G5984GAT_2311_ngat) );
INVXL U_g4665 (.A(G5979GAT_2305_gat), .Y(G5979GAT_2305_ngat) );
INVXL U_g4666 (.A(G5980GAT_2306_gat), .Y(G5980GAT_2306_ngat) );
INVXL U_g4667 (.A(G5975GAT_2307_gat), .Y(G5975GAT_2307_ngat) );
INVXL U_g4668 (.A(G5981GAT_2304_gat), .Y(G5981GAT_2304_ngat) );
INVXL U_g4669 (.A(G732GAT_224_gat), .Y(G732GAT_224_ngat) );
INVXL U_g4670 (.A(G5972GAT_2308_gat), .Y(G5972GAT_2308_ngat) );
INVXL U_g4671 (.A(G5930GAT_2295_gat), .Y(G5930GAT_2295_ngat) );
INVXL U_g4672 (.A(G6030GAT_2313_gat), .Y(G6030GAT_2313_ngat) );
INVXL U_g4673 (.A(G6031GAT_2314_gat), .Y(G6031GAT_2314_ngat) );
INVXL U_g4674 (.A(G6026GAT_2315_gat), .Y(G6026GAT_2315_ngat) );
INVXL U_g4675 (.A(G6023GAT_2316_gat), .Y(G6023GAT_2316_ngat) );
INVXL U_g4676 (.A(G6020GAT_2317_gat), .Y(G6020GAT_2317_ngat) );
INVXL U_g4677 (.A(G6018GAT_2318_gat), .Y(G6018GAT_2318_ngat) );
INVXL U_g4678 (.A(G6019GAT_2321_gat), .Y(G6019GAT_2321_ngat) );
INVXL U_g4679 (.A(G6014GAT_2322_gat), .Y(G6014GAT_2322_ngat) );
INVXL U_g4680 (.A(G6009GAT_2320_gat), .Y(G6009GAT_2320_ngat) );
INVXL U_g4681 (.A(G6010GAT_2323_gat), .Y(G6010GAT_2323_ngat) );
INVXL U_g4682 (.A(G6005GAT_2324_gat), .Y(G6005GAT_2324_ngat) );
INVXL U_g4683 (.A(G6011GAT_2319_gat), .Y(G6011GAT_2319_ngat) );
INVXL U_g4684 (.A(G684GAT_240_gat), .Y(G684GAT_240_ngat) );
INVXL U_g4685 (.A(G6056GAT_2326_gat), .Y(G6056GAT_2326_ngat) );
INVXL U_g4686 (.A(G6057GAT_2327_gat), .Y(G6057GAT_2327_ngat) );
INVXL U_g4687 (.A(G6052GAT_2328_gat), .Y(G6052GAT_2328_ngat) );
INVXL U_g4688 (.A(G6049GAT_2329_gat), .Y(G6049GAT_2329_ngat) );
INVXL U_g4689 (.A(G6046GAT_2330_gat), .Y(G6046GAT_2330_ngat) );
INVXL U_g4690 (.A(G6044GAT_2331_gat), .Y(G6044GAT_2331_ngat) );
INVXL U_g4691 (.A(G6045GAT_2334_gat), .Y(G6045GAT_2334_ngat) );
INVXL U_g4692 (.A(G6040GAT_2335_gat), .Y(G6040GAT_2335_ngat) );
INVXL U_g4693 (.A(G6035GAT_2333_gat), .Y(G6035GAT_2333_ngat) );
INVXL U_g4694 (.A(G6036GAT_2336_gat), .Y(G6036GAT_2336_ngat) );
INVXL U_g4695 (.A(G6037GAT_2332_gat), .Y(G6037GAT_2332_ngat) );
INVXL U_g4696 (.A(G636GAT_256_gat), .Y(G636GAT_256_ngat) );
INVXL U_g4697 (.A(G6080GAT_2338_gat), .Y(G6080GAT_2338_ngat) );
INVXL U_g4698 (.A(G6081GAT_2339_gat), .Y(G6081GAT_2339_ngat) );
INVXL U_g4699 (.A(G6076GAT_2340_gat), .Y(G6076GAT_2340_ngat) );
INVXL U_g4700 (.A(G6073GAT_2341_gat), .Y(G6073GAT_2341_ngat) );
INVXL U_g4701 (.A(G6070GAT_2342_gat), .Y(G6070GAT_2342_ngat) );
INVXL U_g4702 (.A(G6068GAT_2343_gat), .Y(G6068GAT_2343_ngat) );
INVXL U_g4703 (.A(G6069GAT_2345_gat), .Y(G6069GAT_2345_ngat) );
INVXL U_g4704 (.A(G6064GAT_2346_gat), .Y(G6064GAT_2346_ngat) );
INVXL U_g4705 (.A(G6061GAT_2344_gat), .Y(G6061GAT_2344_ngat) );
INVXL U_g4706 (.A(G588GAT_272_gat), .Y(G588GAT_272_ngat) );
INVXL U_g4707 (.A(G6101GAT_2348_gat), .Y(G6101GAT_2348_ngat) );
INVXL U_g4708 (.A(G6102GAT_2349_gat), .Y(G6102GAT_2349_ngat) );
INVXL U_g4709 (.A(G6097GAT_2350_gat), .Y(G6097GAT_2350_ngat) );
INVXL U_g4710 (.A(G6094GAT_2351_gat), .Y(G6094GAT_2351_ngat) );
INVXL U_g4711 (.A(G6091GAT_2352_gat), .Y(G6091GAT_2352_ngat) );
INVXL U_g4712 (.A(G6089GAT_2353_gat), .Y(G6089GAT_2353_ngat) );
INVXL U_g4713 (.A(G6090GAT_2354_gat), .Y(G6090GAT_2354_ngat) );
INVXL U_g4714 (.A(G6085GAT_2355_gat), .Y(G6085GAT_2355_ngat) );
INVXL U_g4715 (.A(G6118GAT_2357_gat), .Y(G6118GAT_2357_ngat) );
INVXL U_g4716 (.A(G6119GAT_2358_gat), .Y(G6119GAT_2358_ngat) );
INVXL U_g4717 (.A(G6114GAT_2359_gat), .Y(G6114GAT_2359_ngat) );
INVXL U_g4718 (.A(G6111GAT_2360_gat), .Y(G6111GAT_2360_ngat) );
INVXL U_g4719 (.A(G6108GAT_2362_gat), .Y(G6108GAT_2362_ngat) );
INVXL U_g4720 (.A(G6106GAT_2361_gat), .Y(G6106GAT_2361_ngat) );
INVXL U_g4721 (.A(G6107GAT_2363_gat), .Y(G6107GAT_2363_ngat) );
INVXL U_g4722 (.A(G6128GAT_2365_gat), .Y(G6128GAT_2365_ngat) );
INVXL U_g4723 (.A(G6129GAT_2366_gat), .Y(G6129GAT_2366_ngat) );
INVXL U_g4724 (.A(G6124GAT_2367_gat), .Y(G6124GAT_2367_ngat) );
INVXL U_g4725 (.A(G6133GAT_2370_gat), .Y(G6133GAT_2370_ngat) );
INVXL U_g4726 (.A(G6134GAT_2371_gat), .Y(G6134GAT_2371_ngat) );
INVXL U_g4727 (.A(G6141GAT_2373_gat), .Y(G6141GAT_2373_ngat) );
INVXL U_g4728 (.A(G6138GAT_2372_gat), .Y(G6138GAT_2372_ngat) );
INVXL U_g4729 (.A(G6135GAT_2369_gat), .Y(G6135GAT_2369_ngat) );
INVXL U_g4730 (.A(G6147GAT_2374_gat), .Y(G6147GAT_2374_ngat) );
INVXL U_g4731 (.A(G6145GAT_2375_gat), .Y(G6145GAT_2375_ngat) );
INVXL U_g4732 (.A(G6146GAT_2376_gat), .Y(G6146GAT_2376_ngat) );
INVXL U_g4733 (.A(G6151GAT_2377_gat), .Y(G6151GAT_2377_ngat) );
INVXL U_g4734 (.A(G6130GAT_2364_gat), .Y(G6130GAT_2364_ngat) );
INVXL U_g4735 (.A(G6157GAT_2379_gat), .Y(G6157GAT_2379_ngat) );
INVXL U_g4736 (.A(G6155GAT_2380_gat), .Y(G6155GAT_2380_ngat) );
INVXL U_g4737 (.A(G6156GAT_2381_gat), .Y(G6156GAT_2381_ngat) );
INVXL U_g4738 (.A(G6161GAT_2382_gat), .Y(G6161GAT_2382_ngat) );
INVXL U_g4739 (.A(G6120GAT_2356_gat), .Y(G6120GAT_2356_ngat) );
INVXL U_g4740 (.A(G6167GAT_2384_gat), .Y(G6167GAT_2384_ngat) );
INVXL U_g4741 (.A(G6165GAT_2385_gat), .Y(G6165GAT_2385_ngat) );
INVXL U_g4742 (.A(G6166GAT_2386_gat), .Y(G6166GAT_2386_ngat) );
INVXL U_g4743 (.A(G6171GAT_2387_gat), .Y(G6171GAT_2387_ngat) );
INVXL U_g4744 (.A(G6103GAT_2347_gat), .Y(G6103GAT_2347_ngat) );
INVXL U_g4745 (.A(G6177GAT_2389_gat), .Y(G6177GAT_2389_ngat) );
INVXL U_g4746 (.A(G6175GAT_2390_gat), .Y(G6175GAT_2390_ngat) );
INVXL U_g4747 (.A(G6176GAT_2391_gat), .Y(G6176GAT_2391_ngat) );
INVXL U_g4748 (.A(G6181GAT_2392_gat), .Y(G6181GAT_2392_ngat) );
INVXL U_g4749 (.A(G6082GAT_2337_gat), .Y(G6082GAT_2337_ngat) );
INVXL U_g4750 (.A(G6187GAT_2394_gat), .Y(G6187GAT_2394_ngat) );
INVXL U_g4751 (.A(G6185GAT_2395_gat), .Y(G6185GAT_2395_ngat) );
INVXL U_g4752 (.A(G6186GAT_2396_gat), .Y(G6186GAT_2396_ngat) );
INVXL U_g4753 (.A(G6191GAT_2397_gat), .Y(G6191GAT_2397_ngat) );
INVXL U_g4754 (.A(G6058GAT_2325_gat), .Y(G6058GAT_2325_ngat) );
INVXL U_g4755 (.A(G6197GAT_2399_gat), .Y(G6197GAT_2399_ngat) );
INVXL U_g4756 (.A(G6195GAT_2400_gat), .Y(G6195GAT_2400_ngat) );
INVXL U_g4757 (.A(G6196GAT_2401_gat), .Y(G6196GAT_2401_ngat) );
INVXL U_g4758 (.A(G6201GAT_2402_gat), .Y(G6201GAT_2402_ngat) );
INVXL U_g4759 (.A(G6032GAT_2312_gat), .Y(G6032GAT_2312_ngat) );
INVXL U_g4760 (.A(G6207GAT_2404_gat), .Y(G6207GAT_2404_ngat) );
INVXL U_g4761 (.A(G6205GAT_2405_gat), .Y(G6205GAT_2405_ngat) );
INVXL U_g4762 (.A(G6206GAT_2406_gat), .Y(G6206GAT_2406_ngat) );
INVXL U_g4763 (.A(G6211GAT_2407_gat), .Y(G6211GAT_2407_ngat) );
INVXL U_g4764 (.A(G6002GAT_2297_gat), .Y(G6002GAT_2297_ngat) );
INVXL U_g4765 (.A(G6217GAT_2409_gat), .Y(G6217GAT_2409_ngat) );
INVXL U_g4766 (.A(G6215GAT_2410_gat), .Y(G6215GAT_2410_ngat) );
INVXL U_g4767 (.A(G6216GAT_2411_gat), .Y(G6216GAT_2411_ngat) );
INVXL U_g4768 (.A(G6221GAT_2412_gat), .Y(G6221GAT_2412_ngat) );
INVXL U_g4769 (.A(G5968GAT_2277_gat), .Y(G5968GAT_2277_ngat) );
INVXL U_g4770 (.A(G6227GAT_2414_gat), .Y(G6227GAT_2414_ngat) );
INVXL U_g4771 (.A(G6225GAT_2415_gat), .Y(G6225GAT_2415_ngat) );
INVXL U_g4772 (.A(G6226GAT_2416_gat), .Y(G6226GAT_2416_ngat) );
INVXL U_g4773 (.A(G6231GAT_2417_gat), .Y(G6231GAT_2417_ngat) );
INVXL U_g4774 (.A(G5925GAT_2258_gat), .Y(G5925GAT_2258_ngat) );
INVXL U_g4775 (.A(G6237GAT_2419_gat), .Y(G6237GAT_2419_ngat) );
INVXL U_g4776 (.A(G6235GAT_2420_gat), .Y(G6235GAT_2420_ngat) );
INVXL U_g4777 (.A(G6236GAT_2421_gat), .Y(G6236GAT_2421_ngat) );
INVXL U_g4778 (.A(G6241GAT_2422_gat), .Y(G6241GAT_2422_ngat) );
INVXL U_g4779 (.A(G5879GAT_2238_gat), .Y(G5879GAT_2238_ngat) );
INVXL U_g4780 (.A(G6247GAT_2424_gat), .Y(G6247GAT_2424_ngat) );
INVXL U_g4781 (.A(G6245GAT_2425_gat), .Y(G6245GAT_2425_ngat) );
INVXL U_g4782 (.A(G6246GAT_2426_gat), .Y(G6246GAT_2426_ngat) );
INVXL U_g4783 (.A(G6251GAT_2427_gat), .Y(G6251GAT_2427_ngat) );
INVXL U_g4784 (.A(G5831GAT_2215_gat), .Y(G5831GAT_2215_ngat) );
INVXL U_g4785 (.A(G6257GAT_2429_gat), .Y(G6257GAT_2429_ngat) );
INVXL U_g4786 (.A(G6255GAT_2430_gat), .Y(G6255GAT_2430_ngat) );
INVXL U_g4787 (.A(G6256GAT_2431_gat), .Y(G6256GAT_2431_ngat) );
INVXL U_g4788 (.A(G6261GAT_2432_gat), .Y(G6261GAT_2432_ngat) );
INVXL U_g4789 (.A(G5782GAT_2192_gat), .Y(G5782GAT_2192_ngat) );
INVXL U_g4790 (.A(G6267GAT_2434_gat), .Y(G6267GAT_2434_ngat) );
INVXL U_g4791 (.A(G6265GAT_2435_gat), .Y(G6265GAT_2435_ngat) );
INVXL U_g4792 (.A(G6266GAT_2436_gat), .Y(G6266GAT_2436_ngat) );
INVXL U_g4793 (.A(G6271GAT_2437_gat), .Y(G6271GAT_2437_ngat) );
INVXL U_g4794 (.A(G5727GAT_2167_gat), .Y(G5727GAT_2167_ngat) );
INVXL U_g4795 (.A(G6277GAT_2439_gat), .Y(G6277GAT_2439_ngat) );
INVXL U_g4796 (.A(G6275GAT_2440_gat), .Y(G6275GAT_2440_ngat) );
INVXL U_g4797 (.A(G6276GAT_2441_gat), .Y(G6276GAT_2441_ngat) );
INVXL U_g4798 (.A(G6281GAT_2442_gat), .Y(G6281GAT_2442_ngat) );
INVXL U_g4799 (.A(G6285GAT_2445_gat), .Y(G6285GAT_2445_ngat) );
INVXL U_g4800 (.A(G6286GAT_2446_gat), .Y(G6286GAT_2446_ngat) );

endmodule
