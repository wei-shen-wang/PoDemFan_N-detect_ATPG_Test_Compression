module C1355 ( G1GAT_0_gat, G8GAT_1_gat, G15GAT_2_gat, G22GAT_3_gat, G29GAT_4_gat, G36GAT_5_gat, G43GAT_6_gat, G50GAT_7_gat, G57GAT_8_gat, G64GAT_9_gat, G71GAT_10_gat, G78GAT_11_gat, G85GAT_12_gat, G92GAT_13_gat, G99GAT_14_gat, G106GAT_15_gat, G113GAT_16_gat, G120GAT_17_gat, G127GAT_18_gat, G134GAT_19_gat, G141GAT_20_gat, G148GAT_21_gat, G155GAT_22_gat, G162GAT_23_gat, G169GAT_24_gat, G176GAT_25_gat, G183GAT_26_gat, G190GAT_27_gat, G197GAT_28_gat, G204GAT_29_gat, G211GAT_30_gat, G218GAT_31_gat, G225GAT_32_gat, G226GAT_33_gat, G227GAT_34_gat, G228GAT_35_gat, G229GAT_36_gat, G230GAT_37_gat, G231GAT_38_gat, G232GAT_39_gat, G233GAT_40_gat, G1324GAT_583_gat, G1325GAT_579_gat, G1326GAT_575_gat, G1327GAT_571_gat, G1328GAT_584_gat, G1329GAT_580_gat, G1330GAT_576_gat, G1331GAT_572_gat, G1332GAT_585_gat, G1333GAT_581_gat, G1334GAT_577_gat, G1335GAT_573_gat, G1336GAT_586_gat, G1337GAT_582_gat, G1338GAT_578_gat, G1339GAT_574_gat, G1340GAT_567_gat, G1341GAT_563_gat, G1342GAT_559_gat, G1343GAT_555_gat, G1344GAT_568_gat, G1345GAT_564_gat, G1346GAT_560_gat, G1347GAT_556_gat, G1348GAT_569_gat, G1349GAT_565_gat, G1350GAT_561_gat, G1351GAT_557_gat, G1352GAT_570_gat, G1353GAT_566_gat, G1354GAT_562_gat, G1355GAT_558_gat);

input G1GAT_0_gat;
input G8GAT_1_gat;
input G15GAT_2_gat;
input G22GAT_3_gat;
input G29GAT_4_gat;
input G36GAT_5_gat;
input G43GAT_6_gat;
input G50GAT_7_gat;
input G57GAT_8_gat;
input G64GAT_9_gat;
input G71GAT_10_gat;
input G78GAT_11_gat;
input G85GAT_12_gat;
input G92GAT_13_gat;
input G99GAT_14_gat;
input G106GAT_15_gat;
input G113GAT_16_gat;
input G120GAT_17_gat;
input G127GAT_18_gat;
input G134GAT_19_gat;
input G141GAT_20_gat;
input G148GAT_21_gat;
input G155GAT_22_gat;
input G162GAT_23_gat;
input G169GAT_24_gat;
input G176GAT_25_gat;
input G183GAT_26_gat;
input G190GAT_27_gat;
input G197GAT_28_gat;
input G204GAT_29_gat;
input G211GAT_30_gat;
input G218GAT_31_gat;
input G225GAT_32_gat;
input G226GAT_33_gat;
input G227GAT_34_gat;
input G228GAT_35_gat;
input G229GAT_36_gat;
input G230GAT_37_gat;
input G231GAT_38_gat;
input G232GAT_39_gat;
input G233GAT_40_gat;

output G1324GAT_583_gat;
output G1325GAT_579_gat;
output G1326GAT_575_gat;
output G1327GAT_571_gat;
output G1328GAT_584_gat;
output G1329GAT_580_gat;
output G1330GAT_576_gat;
output G1331GAT_572_gat;
output G1332GAT_585_gat;
output G1333GAT_581_gat;
output G1334GAT_577_gat;
output G1335GAT_573_gat;
output G1336GAT_586_gat;
output G1337GAT_582_gat;
output G1338GAT_578_gat;
output G1339GAT_574_gat;
output G1340GAT_567_gat;
output G1341GAT_563_gat;
output G1342GAT_559_gat;
output G1343GAT_555_gat;
output G1344GAT_568_gat;
output G1345GAT_564_gat;
output G1346GAT_560_gat;
output G1347GAT_556_gat;
output G1348GAT_569_gat;
output G1349GAT_565_gat;
output G1350GAT_561_gat;
output G1351GAT_557_gat;
output G1352GAT_570_gat;
output G1353GAT_566_gat;
output G1354GAT_562_gat;
output G1355GAT_558_gat;

AND2XL U_g1 (.A(G233GAT_40_gat), .B(G232GAT_39_gat), .Y(G263GAT_41_gat) );
AND2XL U_g2 (.A(G233GAT_40_gat), .B(G231GAT_38_gat), .Y(G260GAT_42_gat) );
AND2XL U_g3 (.A(G233GAT_40_gat), .B(G230GAT_37_gat), .Y(G257GAT_43_gat) );
AND2XL U_g4 (.A(G233GAT_40_gat), .B(G229GAT_36_gat), .Y(G254GAT_44_gat) );
AND2XL U_g5 (.A(G233GAT_40_gat), .B(G228GAT_35_gat), .Y(G251GAT_45_gat) );
AND2XL U_g6 (.A(G233GAT_40_gat), .B(G227GAT_34_gat), .Y(G248GAT_46_gat) );
AND2XL U_g7 (.A(G233GAT_40_gat), .B(G226GAT_33_gat), .Y(G245GAT_47_gat) );
AND2XL U_g8 (.A(G233GAT_40_gat), .B(G225GAT_32_gat), .Y(G242GAT_48_gat) );
AND2XL U_g9 (.A(G218GAT_31_gat), .B(G211GAT_30_gat), .Y(G311GAT_49_gat) );
AND2XL U_g10 (.A(G204GAT_29_gat), .B(G197GAT_28_gat), .Y(G308GAT_50_gat) );
AND2XL U_g11 (.A(G218GAT_31_gat), .B(G190GAT_27_gat), .Y(G359GAT_51_gat) );
AND2XL U_g12 (.A(G211GAT_30_gat), .B(G183GAT_26_gat), .Y(G353GAT_52_gat) );
AND2XL U_g13 (.A(G190GAT_27_gat), .B(G183GAT_26_gat), .Y(G305GAT_53_gat) );
AND2XL U_g14 (.A(G204GAT_29_gat), .B(G176GAT_25_gat), .Y(G347GAT_54_gat) );
AND2XL U_g15 (.A(G197GAT_28_gat), .B(G169GAT_24_gat), .Y(G341GAT_55_gat) );
AND2XL U_g16 (.A(G176GAT_25_gat), .B(G169GAT_24_gat), .Y(G302GAT_56_gat) );
AND2XL U_g17 (.A(G162GAT_23_gat), .B(G155GAT_22_gat), .Y(G299GAT_57_gat) );
AND2XL U_g18 (.A(G148GAT_21_gat), .B(G141GAT_20_gat), .Y(G296GAT_58_gat) );
AND2XL U_g19 (.A(G162GAT_23_gat), .B(G134GAT_19_gat), .Y(G356GAT_59_gat) );
AND2XL U_g20 (.A(G155GAT_22_gat), .B(G127GAT_18_gat), .Y(G350GAT_60_gat) );
AND2XL U_g21 (.A(G134GAT_19_gat), .B(G127GAT_18_gat), .Y(G293GAT_61_gat) );
AND2XL U_g22 (.A(G148GAT_21_gat), .B(G120GAT_17_gat), .Y(G344GAT_62_gat) );
AND2XL U_g23 (.A(G141GAT_20_gat), .B(G113GAT_16_gat), .Y(G338GAT_63_gat) );
AND2XL U_g24 (.A(G120GAT_17_gat), .B(G113GAT_16_gat), .Y(G290GAT_64_gat) );
AND2XL U_g25 (.A(G106GAT_15_gat), .B(G99GAT_14_gat), .Y(G287GAT_65_gat) );
AND2XL U_g26 (.A(G92GAT_13_gat), .B(G85GAT_12_gat), .Y(G284GAT_66_gat) );
AND2XL U_g27 (.A(G106GAT_15_gat), .B(G78GAT_11_gat), .Y(G335GAT_67_gat) );
AND2XL U_g28 (.A(G99GAT_14_gat), .B(G71GAT_10_gat), .Y(G329GAT_68_gat) );
AND2XL U_g29 (.A(G78GAT_11_gat), .B(G71GAT_10_gat), .Y(G281GAT_69_gat) );
AND2XL U_g30 (.A(G92GAT_13_gat), .B(G64GAT_9_gat), .Y(G323GAT_70_gat) );
AND2XL U_g31 (.A(G85GAT_12_gat), .B(G57GAT_8_gat), .Y(G317GAT_71_gat) );
AND2XL U_g32 (.A(G64GAT_9_gat), .B(G57GAT_8_gat), .Y(G278GAT_72_gat) );
AND2XL U_g33 (.A(G50GAT_7_gat), .B(G43GAT_6_gat), .Y(G275GAT_73_gat) );
AND2XL U_g34 (.A(G36GAT_5_gat), .B(G29GAT_4_gat), .Y(G272GAT_74_gat) );
AND2XL U_g35 (.A(G50GAT_7_gat), .B(G22GAT_3_gat), .Y(G332GAT_75_gat) );
AND2XL U_g36 (.A(G43GAT_6_gat), .B(G15GAT_2_gat), .Y(G326GAT_76_gat) );
AND2XL U_g37 (.A(G22GAT_3_gat), .B(G15GAT_2_gat), .Y(G269GAT_77_gat) );
AND2XL U_g38 (.A(G36GAT_5_gat), .B(G8GAT_1_gat), .Y(G320GAT_78_gat) );
AND2XL U_g39 (.A(G29GAT_4_gat), .B(G1GAT_0_gat), .Y(G314GAT_79_gat) );
AND2XL U_g40 (.A(G8GAT_1_gat), .B(G1GAT_0_gat), .Y(G266GAT_80_gat) );
AND2XL U_g41 (.A(G359GAT_51_gat), .B(G218GAT_31_gat), .Y(G425GAT_81_gat) );
AND2XL U_g42 (.A(G311GAT_49_gat), .B(G218GAT_31_gat), .Y(G393GAT_82_gat) );
AND2XL U_g43 (.A(G353GAT_52_gat), .B(G211GAT_30_gat), .Y(G421GAT_83_gat) );
AND2XL U_g44 (.A(G311GAT_49_gat), .B(G211GAT_30_gat), .Y(G392GAT_84_gat) );
AND2XL U_g45 (.A(G347GAT_54_gat), .B(G204GAT_29_gat), .Y(G417GAT_85_gat) );
AND2XL U_g46 (.A(G308GAT_50_gat), .B(G204GAT_29_gat), .Y(G391GAT_86_gat) );
AND2XL U_g47 (.A(G341GAT_55_gat), .B(G197GAT_28_gat), .Y(G413GAT_87_gat) );
AND2XL U_g48 (.A(G308GAT_50_gat), .B(G197GAT_28_gat), .Y(G390GAT_88_gat) );
AND2XL U_g49 (.A(G359GAT_51_gat), .B(G190GAT_27_gat), .Y(G424GAT_89_gat) );
AND2XL U_g50 (.A(G305GAT_53_gat), .B(G190GAT_27_gat), .Y(G389GAT_90_gat) );
AND2XL U_g51 (.A(G353GAT_52_gat), .B(G183GAT_26_gat), .Y(G420GAT_91_gat) );
AND2XL U_g52 (.A(G305GAT_53_gat), .B(G183GAT_26_gat), .Y(G388GAT_92_gat) );
AND2XL U_g53 (.A(G347GAT_54_gat), .B(G176GAT_25_gat), .Y(G416GAT_93_gat) );
AND2XL U_g54 (.A(G302GAT_56_gat), .B(G176GAT_25_gat), .Y(G387GAT_94_gat) );
AND2XL U_g55 (.A(G341GAT_55_gat), .B(G169GAT_24_gat), .Y(G412GAT_95_gat) );
AND2XL U_g56 (.A(G302GAT_56_gat), .B(G169GAT_24_gat), .Y(G386GAT_96_gat) );
AND2XL U_g57 (.A(G356GAT_59_gat), .B(G162GAT_23_gat), .Y(G423GAT_97_gat) );
AND2XL U_g58 (.A(G299GAT_57_gat), .B(G162GAT_23_gat), .Y(G385GAT_98_gat) );
AND2XL U_g59 (.A(G350GAT_60_gat), .B(G155GAT_22_gat), .Y(G419GAT_99_gat) );
AND2XL U_g60 (.A(G299GAT_57_gat), .B(G155GAT_22_gat), .Y(G384GAT_100_gat) );
AND2XL U_g61 (.A(G344GAT_62_gat), .B(G148GAT_21_gat), .Y(G415GAT_101_gat) );
AND2XL U_g62 (.A(G296GAT_58_gat), .B(G148GAT_21_gat), .Y(G383GAT_102_gat) );
AND2XL U_g63 (.A(G338GAT_63_gat), .B(G141GAT_20_gat), .Y(G411GAT_103_gat) );
AND2XL U_g64 (.A(G296GAT_58_gat), .B(G141GAT_20_gat), .Y(G382GAT_104_gat) );
AND2XL U_g65 (.A(G356GAT_59_gat), .B(G134GAT_19_gat), .Y(G422GAT_105_gat) );
AND2XL U_g66 (.A(G293GAT_61_gat), .B(G134GAT_19_gat), .Y(G381GAT_106_gat) );
AND2XL U_g67 (.A(G350GAT_60_gat), .B(G127GAT_18_gat), .Y(G418GAT_107_gat) );
AND2XL U_g68 (.A(G293GAT_61_gat), .B(G127GAT_18_gat), .Y(G380GAT_108_gat) );
AND2XL U_g69 (.A(G344GAT_62_gat), .B(G120GAT_17_gat), .Y(G414GAT_109_gat) );
AND2XL U_g70 (.A(G290GAT_64_gat), .B(G120GAT_17_gat), .Y(G379GAT_110_gat) );
AND2XL U_g71 (.A(G338GAT_63_gat), .B(G113GAT_16_gat), .Y(G410GAT_111_gat) );
AND2XL U_g72 (.A(G290GAT_64_gat), .B(G113GAT_16_gat), .Y(G378GAT_112_gat) );
AND2XL U_g73 (.A(G335GAT_67_gat), .B(G106GAT_15_gat), .Y(G409GAT_113_gat) );
AND2XL U_g74 (.A(G287GAT_65_gat), .B(G106GAT_15_gat), .Y(G377GAT_114_gat) );
AND2XL U_g75 (.A(G329GAT_68_gat), .B(G99GAT_14_gat), .Y(G405GAT_115_gat) );
AND2XL U_g76 (.A(G287GAT_65_gat), .B(G99GAT_14_gat), .Y(G376GAT_116_gat) );
AND2XL U_g77 (.A(G323GAT_70_gat), .B(G92GAT_13_gat), .Y(G401GAT_117_gat) );
AND2XL U_g78 (.A(G284GAT_66_gat), .B(G92GAT_13_gat), .Y(G375GAT_118_gat) );
AND2XL U_g79 (.A(G317GAT_71_gat), .B(G85GAT_12_gat), .Y(G397GAT_119_gat) );
AND2XL U_g80 (.A(G284GAT_66_gat), .B(G85GAT_12_gat), .Y(G374GAT_120_gat) );
AND2XL U_g81 (.A(G335GAT_67_gat), .B(G78GAT_11_gat), .Y(G408GAT_121_gat) );
AND2XL U_g82 (.A(G281GAT_69_gat), .B(G78GAT_11_gat), .Y(G373GAT_122_gat) );
AND2XL U_g83 (.A(G329GAT_68_gat), .B(G71GAT_10_gat), .Y(G404GAT_123_gat) );
AND2XL U_g84 (.A(G281GAT_69_gat), .B(G71GAT_10_gat), .Y(G372GAT_124_gat) );
AND2XL U_g85 (.A(G323GAT_70_gat), .B(G64GAT_9_gat), .Y(G400GAT_125_gat) );
AND2XL U_g86 (.A(G278GAT_72_gat), .B(G64GAT_9_gat), .Y(G371GAT_126_gat) );
AND2XL U_g87 (.A(G317GAT_71_gat), .B(G57GAT_8_gat), .Y(G396GAT_127_gat) );
AND2XL U_g88 (.A(G278GAT_72_gat), .B(G57GAT_8_gat), .Y(G370GAT_128_gat) );
AND2XL U_g89 (.A(G332GAT_75_gat), .B(G50GAT_7_gat), .Y(G407GAT_129_gat) );
AND2XL U_g90 (.A(G275GAT_73_gat), .B(G50GAT_7_gat), .Y(G369GAT_130_gat) );
AND2XL U_g91 (.A(G326GAT_76_gat), .B(G43GAT_6_gat), .Y(G403GAT_131_gat) );
AND2XL U_g92 (.A(G275GAT_73_gat), .B(G43GAT_6_gat), .Y(G368GAT_132_gat) );
AND2XL U_g93 (.A(G320GAT_78_gat), .B(G36GAT_5_gat), .Y(G399GAT_133_gat) );
AND2XL U_g94 (.A(G272GAT_74_gat), .B(G36GAT_5_gat), .Y(G367GAT_134_gat) );
AND2XL U_g95 (.A(G314GAT_79_gat), .B(G29GAT_4_gat), .Y(G395GAT_135_gat) );
AND2XL U_g96 (.A(G272GAT_74_gat), .B(G29GAT_4_gat), .Y(G366GAT_136_gat) );
AND2XL U_g97 (.A(G332GAT_75_gat), .B(G22GAT_3_gat), .Y(G406GAT_137_gat) );
AND2XL U_g98 (.A(G269GAT_77_gat), .B(G22GAT_3_gat), .Y(G365GAT_138_gat) );
AND2XL U_g99 (.A(G326GAT_76_gat), .B(G15GAT_2_gat), .Y(G402GAT_139_gat) );
AND2XL U_g100 (.A(G269GAT_77_gat), .B(G15GAT_2_gat), .Y(G364GAT_140_gat) );
AND2XL U_g101 (.A(G320GAT_78_gat), .B(G8GAT_1_gat), .Y(G398GAT_141_gat) );
AND2XL U_g102 (.A(G266GAT_80_gat), .B(G8GAT_1_gat), .Y(G363GAT_142_gat) );
AND2XL U_g103 (.A(G314GAT_79_gat), .B(G1GAT_0_gat), .Y(G394GAT_143_gat) );
AND2XL U_g104 (.A(G266GAT_80_gat), .B(G1GAT_0_gat), .Y(G362GAT_144_gat) );
AND2XL U_g105 (.A(G425GAT_81_gat), .B(G424GAT_89_gat), .Y(G519GAT_145_gat) );
AND2XL U_g106 (.A(G393GAT_82_gat), .B(G392GAT_84_gat), .Y(G471GAT_146_gat) );
AND2XL U_g107 (.A(G421GAT_83_gat), .B(G420GAT_91_gat), .Y(G513GAT_147_gat) );
AND2XL U_g108 (.A(G417GAT_85_gat), .B(G416GAT_93_gat), .Y(G507GAT_148_gat) );
AND2XL U_g109 (.A(G391GAT_86_gat), .B(G390GAT_88_gat), .Y(G468GAT_149_gat) );
AND2XL U_g110 (.A(G413GAT_87_gat), .B(G412GAT_95_gat), .Y(G501GAT_150_gat) );
AND2XL U_g111 (.A(G389GAT_90_gat), .B(G388GAT_92_gat), .Y(G465GAT_151_gat) );
AND2XL U_g112 (.A(G387GAT_94_gat), .B(G386GAT_96_gat), .Y(G462GAT_152_gat) );
AND2XL U_g113 (.A(G423GAT_97_gat), .B(G422GAT_105_gat), .Y(G516GAT_153_gat) );
AND2XL U_g114 (.A(G385GAT_98_gat), .B(G384GAT_100_gat), .Y(G459GAT_154_gat) );
AND2XL U_g115 (.A(G419GAT_99_gat), .B(G418GAT_107_gat), .Y(G510GAT_155_gat) );
AND2XL U_g116 (.A(G415GAT_101_gat), .B(G414GAT_109_gat), .Y(G504GAT_156_gat) );
AND2XL U_g117 (.A(G383GAT_102_gat), .B(G382GAT_104_gat), .Y(G456GAT_157_gat) );
AND2XL U_g118 (.A(G411GAT_103_gat), .B(G410GAT_111_gat), .Y(G498GAT_158_gat) );
AND2XL U_g119 (.A(G381GAT_106_gat), .B(G380GAT_108_gat), .Y(G453GAT_159_gat) );
AND2XL U_g120 (.A(G379GAT_110_gat), .B(G378GAT_112_gat), .Y(G450GAT_160_gat) );
AND2XL U_g121 (.A(G409GAT_113_gat), .B(G408GAT_121_gat), .Y(G495GAT_161_gat) );
AND2XL U_g122 (.A(G377GAT_114_gat), .B(G376GAT_116_gat), .Y(G447GAT_162_gat) );
AND2XL U_g123 (.A(G405GAT_115_gat), .B(G404GAT_123_gat), .Y(G489GAT_163_gat) );
AND2XL U_g124 (.A(G401GAT_117_gat), .B(G400GAT_125_gat), .Y(G483GAT_164_gat) );
AND2XL U_g125 (.A(G375GAT_118_gat), .B(G374GAT_120_gat), .Y(G444GAT_165_gat) );
AND2XL U_g126 (.A(G397GAT_119_gat), .B(G396GAT_127_gat), .Y(G477GAT_166_gat) );
AND2XL U_g127 (.A(G373GAT_122_gat), .B(G372GAT_124_gat), .Y(G441GAT_167_gat) );
AND2XL U_g128 (.A(G371GAT_126_gat), .B(G370GAT_128_gat), .Y(G438GAT_168_gat) );
AND2XL U_g129 (.A(G407GAT_129_gat), .B(G406GAT_137_gat), .Y(G492GAT_169_gat) );
AND2XL U_g130 (.A(G369GAT_130_gat), .B(G368GAT_132_gat), .Y(G435GAT_170_gat) );
AND2XL U_g131 (.A(G403GAT_131_gat), .B(G402GAT_139_gat), .Y(G486GAT_171_gat) );
AND2XL U_g132 (.A(G399GAT_133_gat), .B(G398GAT_141_gat), .Y(G480GAT_172_gat) );
AND2XL U_g133 (.A(G367GAT_134_gat), .B(G366GAT_136_gat), .Y(G432GAT_173_gat) );
AND2XL U_g134 (.A(G395GAT_135_gat), .B(G394GAT_143_gat), .Y(G474GAT_174_gat) );
AND2XL U_g135 (.A(G365GAT_138_gat), .B(G364GAT_140_gat), .Y(G429GAT_175_gat) );
AND2XL U_g136 (.A(G363GAT_142_gat), .B(G362GAT_144_gat), .Y(G426GAT_176_gat) );
AND2XL U_g137 (.A(G519GAT_145_gat), .B(G516GAT_153_gat), .Y(G567GAT_177_gat) );
AND2XL U_g138 (.A(G471GAT_146_gat), .B(G468GAT_149_gat), .Y(G543GAT_178_gat) );
AND2XL U_g139 (.A(G513GAT_147_gat), .B(G510GAT_155_gat), .Y(G564GAT_179_gat) );
AND2XL U_g140 (.A(G507GAT_148_gat), .B(G504GAT_156_gat), .Y(G561GAT_180_gat) );
AND2XL U_g141 (.A(G501GAT_150_gat), .B(G498GAT_158_gat), .Y(G558GAT_181_gat) );
AND2XL U_g142 (.A(G465GAT_151_gat), .B(G462GAT_152_gat), .Y(G540GAT_182_gat) );
AND2XL U_g143 (.A(G459GAT_154_gat), .B(G456GAT_157_gat), .Y(G537GAT_183_gat) );
AND2XL U_g144 (.A(G453GAT_159_gat), .B(G450GAT_160_gat), .Y(G534GAT_184_gat) );
AND2XL U_g145 (.A(G495GAT_161_gat), .B(G492GAT_169_gat), .Y(G555GAT_185_gat) );
AND2XL U_g146 (.A(G447GAT_162_gat), .B(G444GAT_165_gat), .Y(G531GAT_186_gat) );
AND2XL U_g147 (.A(G489GAT_163_gat), .B(G486GAT_171_gat), .Y(G552GAT_187_gat) );
AND2XL U_g148 (.A(G483GAT_164_gat), .B(G480GAT_172_gat), .Y(G549GAT_188_gat) );
AND2XL U_g149 (.A(G477GAT_166_gat), .B(G474GAT_174_gat), .Y(G546GAT_189_gat) );
AND2XL U_g150 (.A(G441GAT_167_gat), .B(G438GAT_168_gat), .Y(G528GAT_190_gat) );
AND2XL U_g151 (.A(G435GAT_170_gat), .B(G432GAT_173_gat), .Y(G525GAT_191_gat) );
AND2XL U_g152 (.A(G429GAT_175_gat), .B(G426GAT_176_gat), .Y(G522GAT_192_gat) );
AND2XL U_g153 (.A(G567GAT_177_gat), .B(G519GAT_145_gat), .Y(G601GAT_193_gat) );
AND2XL U_g154 (.A(G543GAT_178_gat), .B(G471GAT_146_gat), .Y(G585GAT_194_gat) );
AND2XL U_g155 (.A(G564GAT_179_gat), .B(G513GAT_147_gat), .Y(G599GAT_195_gat) );
AND2XL U_g156 (.A(G561GAT_180_gat), .B(G507GAT_148_gat), .Y(G597GAT_196_gat) );
AND2XL U_g157 (.A(G543GAT_178_gat), .B(G468GAT_149_gat), .Y(G584GAT_197_gat) );
AND2XL U_g158 (.A(G558GAT_181_gat), .B(G501GAT_150_gat), .Y(G595GAT_198_gat) );
AND2XL U_g159 (.A(G540GAT_182_gat), .B(G465GAT_151_gat), .Y(G583GAT_199_gat) );
AND2XL U_g160 (.A(G540GAT_182_gat), .B(G462GAT_152_gat), .Y(G582GAT_200_gat) );
AND2XL U_g161 (.A(G567GAT_177_gat), .B(G516GAT_153_gat), .Y(G600GAT_201_gat) );
AND2XL U_g162 (.A(G537GAT_183_gat), .B(G459GAT_154_gat), .Y(G581GAT_202_gat) );
AND2XL U_g163 (.A(G564GAT_179_gat), .B(G510GAT_155_gat), .Y(G598GAT_203_gat) );
AND2XL U_g164 (.A(G561GAT_180_gat), .B(G504GAT_156_gat), .Y(G596GAT_204_gat) );
AND2XL U_g165 (.A(G537GAT_183_gat), .B(G456GAT_157_gat), .Y(G580GAT_205_gat) );
AND2XL U_g166 (.A(G558GAT_181_gat), .B(G498GAT_158_gat), .Y(G594GAT_206_gat) );
AND2XL U_g167 (.A(G534GAT_184_gat), .B(G453GAT_159_gat), .Y(G579GAT_207_gat) );
AND2XL U_g168 (.A(G534GAT_184_gat), .B(G450GAT_160_gat), .Y(G578GAT_208_gat) );
AND2XL U_g169 (.A(G555GAT_185_gat), .B(G495GAT_161_gat), .Y(G593GAT_209_gat) );
AND2XL U_g170 (.A(G531GAT_186_gat), .B(G447GAT_162_gat), .Y(G577GAT_210_gat) );
AND2XL U_g171 (.A(G552GAT_187_gat), .B(G489GAT_163_gat), .Y(G591GAT_211_gat) );
AND2XL U_g172 (.A(G549GAT_188_gat), .B(G483GAT_164_gat), .Y(G589GAT_212_gat) );
AND2XL U_g173 (.A(G531GAT_186_gat), .B(G444GAT_165_gat), .Y(G576GAT_213_gat) );
AND2XL U_g174 (.A(G546GAT_189_gat), .B(G477GAT_166_gat), .Y(G587GAT_214_gat) );
AND2XL U_g175 (.A(G528GAT_190_gat), .B(G441GAT_167_gat), .Y(G575GAT_215_gat) );
AND2XL U_g176 (.A(G528GAT_190_gat), .B(G438GAT_168_gat), .Y(G574GAT_216_gat) );
AND2XL U_g177 (.A(G555GAT_185_gat), .B(G492GAT_169_gat), .Y(G592GAT_217_gat) );
AND2XL U_g178 (.A(G525GAT_191_gat), .B(G435GAT_170_gat), .Y(G573GAT_218_gat) );
AND2XL U_g179 (.A(G552GAT_187_gat), .B(G486GAT_171_gat), .Y(G590GAT_219_gat) );
AND2XL U_g180 (.A(G549GAT_188_gat), .B(G480GAT_172_gat), .Y(G588GAT_220_gat) );
AND2XL U_g181 (.A(G525GAT_191_gat), .B(G432GAT_173_gat), .Y(G572GAT_221_gat) );
AND2XL U_g182 (.A(G546GAT_189_gat), .B(G474GAT_174_gat), .Y(G586GAT_222_gat) );
AND2XL U_g183 (.A(G522GAT_192_gat), .B(G429GAT_175_gat), .Y(G571GAT_223_gat) );
AND2XL U_g184 (.A(G522GAT_192_gat), .B(G426GAT_176_gat), .Y(G570GAT_224_gat) );
AND2XL U_g185 (.A(G601GAT_193_gat), .B(G600GAT_201_gat), .Y(G663GAT_225_gat) );
AND2XL U_g186 (.A(G585GAT_194_gat), .B(G584GAT_197_gat), .Y(G637GAT_226_gat) );
AND2XL U_g187 (.A(G599GAT_195_gat), .B(G598GAT_203_gat), .Y(G660GAT_227_gat) );
AND2XL U_g188 (.A(G597GAT_196_gat), .B(G596GAT_204_gat), .Y(G657GAT_228_gat) );
AND2XL U_g189 (.A(G595GAT_198_gat), .B(G594GAT_206_gat), .Y(G654GAT_229_gat) );
AND2XL U_g190 (.A(G583GAT_199_gat), .B(G582GAT_200_gat), .Y(G632GAT_230_gat) );
AND2XL U_g191 (.A(G581GAT_202_gat), .B(G580GAT_205_gat), .Y(G627GAT_231_gat) );
AND2XL U_g192 (.A(G579GAT_207_gat), .B(G578GAT_208_gat), .Y(G622GAT_232_gat) );
AND2XL U_g193 (.A(G593GAT_209_gat), .B(G592GAT_217_gat), .Y(G651GAT_233_gat) );
AND2XL U_g194 (.A(G577GAT_210_gat), .B(G576GAT_213_gat), .Y(G617GAT_234_gat) );
AND2XL U_g195 (.A(G591GAT_211_gat), .B(G590GAT_219_gat), .Y(G648GAT_235_gat) );
AND2XL U_g196 (.A(G589GAT_212_gat), .B(G588GAT_220_gat), .Y(G645GAT_236_gat) );
AND2XL U_g197 (.A(G587GAT_214_gat), .B(G586GAT_222_gat), .Y(G642GAT_237_gat) );
AND2XL U_g198 (.A(G575GAT_215_gat), .B(G574GAT_216_gat), .Y(G612GAT_238_gat) );
AND2XL U_g199 (.A(G573GAT_218_gat), .B(G572GAT_221_gat), .Y(G607GAT_239_gat) );
AND2XL U_g200 (.A(G571GAT_223_gat), .B(G570GAT_224_gat), .Y(G602GAT_240_gat) );
AND2XL U_g201 (.A(G637GAT_226_gat), .B(G632GAT_230_gat), .Y(G681GAT_241_gat) );
AND2XL U_g202 (.A(G637GAT_226_gat), .B(G627GAT_231_gat), .Y(G687GAT_242_gat) );
AND2XL U_g203 (.A(G632GAT_230_gat), .B(G622GAT_232_gat), .Y(G684GAT_243_gat) );
AND2XL U_g204 (.A(G627GAT_231_gat), .B(G622GAT_232_gat), .Y(G678GAT_244_gat) );
AND2XL U_g205 (.A(G617GAT_234_gat), .B(G612GAT_238_gat), .Y(G669GAT_245_gat) );
AND2XL U_g206 (.A(G617GAT_234_gat), .B(G607GAT_239_gat), .Y(G675GAT_246_gat) );
AND2XL U_g207 (.A(G612GAT_238_gat), .B(G602GAT_240_gat), .Y(G672GAT_247_gat) );
AND2XL U_g208 (.A(G607GAT_239_gat), .B(G602GAT_240_gat), .Y(G666GAT_248_gat) );
AND2XL U_g209 (.A(G681GAT_241_gat), .B(G637GAT_226_gat), .Y(G701GAT_249_gat) );
AND2XL U_g210 (.A(G687GAT_242_gat), .B(G637GAT_226_gat), .Y(G705GAT_250_gat) );
AND2XL U_g211 (.A(G681GAT_241_gat), .B(G632GAT_230_gat), .Y(G700GAT_251_gat) );
AND2XL U_g212 (.A(G684GAT_243_gat), .B(G632GAT_230_gat), .Y(G703GAT_252_gat) );
AND2XL U_g213 (.A(G678GAT_244_gat), .B(G627GAT_231_gat), .Y(G699GAT_253_gat) );
AND2XL U_g214 (.A(G687GAT_242_gat), .B(G627GAT_231_gat), .Y(G704GAT_254_gat) );
AND2XL U_g215 (.A(G678GAT_244_gat), .B(G622GAT_232_gat), .Y(G698GAT_255_gat) );
AND2XL U_g216 (.A(G684GAT_243_gat), .B(G622GAT_232_gat), .Y(G702GAT_256_gat) );
AND2XL U_g217 (.A(G669GAT_245_gat), .B(G617GAT_234_gat), .Y(G693GAT_257_gat) );
AND2XL U_g218 (.A(G675GAT_246_gat), .B(G617GAT_234_gat), .Y(G697GAT_258_gat) );
AND2XL U_g219 (.A(G669GAT_245_gat), .B(G612GAT_238_gat), .Y(G692GAT_259_gat) );
AND2XL U_g220 (.A(G672GAT_247_gat), .B(G612GAT_238_gat), .Y(G695GAT_260_gat) );
AND2XL U_g221 (.A(G666GAT_248_gat), .B(G607GAT_239_gat), .Y(G691GAT_261_gat) );
AND2XL U_g222 (.A(G675GAT_246_gat), .B(G607GAT_239_gat), .Y(G696GAT_262_gat) );
AND2XL U_g223 (.A(G666GAT_248_gat), .B(G602GAT_240_gat), .Y(G690GAT_263_gat) );
AND2XL U_g224 (.A(G672GAT_247_gat), .B(G602GAT_240_gat), .Y(G694GAT_264_gat) );
AND2XL U_g225 (.A(G701GAT_249_gat), .B(G700GAT_251_gat), .Y(G721GAT_265_gat) );
AND2XL U_g226 (.A(G705GAT_250_gat), .B(G704GAT_254_gat), .Y(G727GAT_266_gat) );
AND2XL U_g227 (.A(G703GAT_252_gat), .B(G702GAT_256_gat), .Y(G724GAT_267_gat) );
AND2XL U_g228 (.A(G699GAT_253_gat), .B(G698GAT_255_gat), .Y(G718GAT_268_gat) );
AND2XL U_g229 (.A(G693GAT_257_gat), .B(G692GAT_259_gat), .Y(G709GAT_269_gat) );
AND2XL U_g230 (.A(G697GAT_258_gat), .B(G696GAT_262_gat), .Y(G715GAT_270_gat) );
AND2XL U_g231 (.A(G695GAT_260_gat), .B(G694GAT_264_gat), .Y(G712GAT_271_gat) );
AND2XL U_g232 (.A(G691GAT_261_gat), .B(G690GAT_263_gat), .Y(G706GAT_272_gat) );
AND2XL U_g233 (.A(G715GAT_270_gat), .B(G263GAT_41_gat), .Y(G751GAT_273_gat) );
AND2XL U_g234 (.A(G712GAT_271_gat), .B(G260GAT_42_gat), .Y(G748GAT_274_gat) );
AND2XL U_g235 (.A(G709GAT_269_gat), .B(G257GAT_43_gat), .Y(G745GAT_275_gat) );
AND2XL U_g236 (.A(G706GAT_272_gat), .B(G254GAT_44_gat), .Y(G742GAT_276_gat) );
AND2XL U_g237 (.A(G727GAT_266_gat), .B(G251GAT_45_gat), .Y(G739GAT_277_gat) );
AND2XL U_g238 (.A(G724GAT_267_gat), .B(G248GAT_46_gat), .Y(G736GAT_278_gat) );
AND2XL U_g239 (.A(G721GAT_265_gat), .B(G245GAT_47_gat), .Y(G733GAT_279_gat) );
AND2XL U_g240 (.A(G718GAT_268_gat), .B(G242GAT_48_gat), .Y(G730GAT_280_gat) );
AND2XL U_g241 (.A(G751GAT_273_gat), .B(G263GAT_41_gat), .Y(G768GAT_281_gat) );
AND2XL U_g242 (.A(G748GAT_274_gat), .B(G260GAT_42_gat), .Y(G766GAT_282_gat) );
AND2XL U_g243 (.A(G745GAT_275_gat), .B(G257GAT_43_gat), .Y(G764GAT_283_gat) );
AND2XL U_g244 (.A(G742GAT_276_gat), .B(G254GAT_44_gat), .Y(G762GAT_284_gat) );
AND2XL U_g245 (.A(G739GAT_277_gat), .B(G251GAT_45_gat), .Y(G760GAT_285_gat) );
AND2XL U_g246 (.A(G736GAT_278_gat), .B(G248GAT_46_gat), .Y(G758GAT_286_gat) );
AND2XL U_g247 (.A(G733GAT_279_gat), .B(G245GAT_47_gat), .Y(G756GAT_287_gat) );
AND2XL U_g248 (.A(G730GAT_280_gat), .B(G242GAT_48_gat), .Y(G754GAT_288_gat) );
AND2XL U_g249 (.A(G733GAT_279_gat), .B(G721GAT_265_gat), .Y(G757GAT_289_gat) );
AND2XL U_g250 (.A(G739GAT_277_gat), .B(G727GAT_266_gat), .Y(G761GAT_290_gat) );
AND2XL U_g251 (.A(G736GAT_278_gat), .B(G724GAT_267_gat), .Y(G759GAT_291_gat) );
AND2XL U_g252 (.A(G730GAT_280_gat), .B(G718GAT_268_gat), .Y(G755GAT_292_gat) );
AND2XL U_g253 (.A(G745GAT_275_gat), .B(G709GAT_269_gat), .Y(G765GAT_293_gat) );
AND2XL U_g254 (.A(G751GAT_273_gat), .B(G715GAT_270_gat), .Y(G769GAT_294_gat) );
AND2XL U_g255 (.A(G748GAT_274_gat), .B(G712GAT_271_gat), .Y(G767GAT_295_gat) );
AND2XL U_g256 (.A(G742GAT_276_gat), .B(G706GAT_272_gat), .Y(G763GAT_296_gat) );
AND2XL U_g257 (.A(G769GAT_294_gat), .B(G768GAT_281_gat), .Y(G791GAT_297_gat) );
AND2XL U_g258 (.A(G767GAT_295_gat), .B(G766GAT_282_gat), .Y(G788GAT_298_gat) );
AND2XL U_g259 (.A(G765GAT_293_gat), .B(G764GAT_283_gat), .Y(G785GAT_299_gat) );
AND2XL U_g260 (.A(G763GAT_296_gat), .B(G762GAT_284_gat), .Y(G782GAT_300_gat) );
AND2XL U_g261 (.A(G761GAT_290_gat), .B(G760GAT_285_gat), .Y(G779GAT_301_gat) );
AND2XL U_g262 (.A(G759GAT_291_gat), .B(G758GAT_286_gat), .Y(G776GAT_302_gat) );
AND2XL U_g263 (.A(G757GAT_289_gat), .B(G756GAT_287_gat), .Y(G773GAT_303_gat) );
AND2XL U_g264 (.A(G755GAT_292_gat), .B(G754GAT_288_gat), .Y(G770GAT_304_gat) );
AND2XL U_g265 (.A(G791GAT_297_gat), .B(G663GAT_225_gat), .Y(G815GAT_305_gat) );
AND2XL U_g266 (.A(G788GAT_298_gat), .B(G660GAT_227_gat), .Y(G812GAT_306_gat) );
AND2XL U_g267 (.A(G785GAT_299_gat), .B(G657GAT_228_gat), .Y(G809GAT_307_gat) );
AND2XL U_g268 (.A(G782GAT_300_gat), .B(G654GAT_229_gat), .Y(G806GAT_308_gat) );
AND2XL U_g269 (.A(G779GAT_301_gat), .B(G651GAT_233_gat), .Y(G803GAT_309_gat) );
AND2XL U_g270 (.A(G776GAT_302_gat), .B(G648GAT_235_gat), .Y(G800GAT_310_gat) );
AND2XL U_g271 (.A(G773GAT_303_gat), .B(G645GAT_236_gat), .Y(G797GAT_311_gat) );
AND2XL U_g272 (.A(G770GAT_304_gat), .B(G642GAT_237_gat), .Y(G794GAT_312_gat) );
AND2XL U_g273 (.A(G815GAT_305_gat), .B(G791GAT_297_gat), .Y(G833GAT_313_gat) );
AND2XL U_g274 (.A(G812GAT_306_gat), .B(G788GAT_298_gat), .Y(G831GAT_314_gat) );
AND2XL U_g275 (.A(G809GAT_307_gat), .B(G785GAT_299_gat), .Y(G829GAT_315_gat) );
AND2XL U_g276 (.A(G806GAT_308_gat), .B(G782GAT_300_gat), .Y(G827GAT_316_gat) );
AND2XL U_g277 (.A(G803GAT_309_gat), .B(G779GAT_301_gat), .Y(G825GAT_317_gat) );
AND2XL U_g278 (.A(G800GAT_310_gat), .B(G776GAT_302_gat), .Y(G823GAT_318_gat) );
AND2XL U_g279 (.A(G797GAT_311_gat), .B(G773GAT_303_gat), .Y(G821GAT_319_gat) );
AND2XL U_g280 (.A(G794GAT_312_gat), .B(G770GAT_304_gat), .Y(G819GAT_320_gat) );
AND2XL U_g281 (.A(G815GAT_305_gat), .B(G663GAT_225_gat), .Y(G832GAT_321_gat) );
AND2XL U_g282 (.A(G812GAT_306_gat), .B(G660GAT_227_gat), .Y(G830GAT_322_gat) );
AND2XL U_g283 (.A(G809GAT_307_gat), .B(G657GAT_228_gat), .Y(G828GAT_323_gat) );
AND2XL U_g284 (.A(G806GAT_308_gat), .B(G654GAT_229_gat), .Y(G826GAT_324_gat) );
AND2XL U_g285 (.A(G803GAT_309_gat), .B(G651GAT_233_gat), .Y(G824GAT_325_gat) );
AND2XL U_g286 (.A(G800GAT_310_gat), .B(G648GAT_235_gat), .Y(G822GAT_326_gat) );
AND2XL U_g287 (.A(G797GAT_311_gat), .B(G645GAT_236_gat), .Y(G820GAT_327_gat) );
AND2XL U_g288 (.A(G794GAT_312_gat), .B(G642GAT_237_gat), .Y(G818GAT_328_gat) );
AND2XL U_g289 (.A(G833GAT_313_gat), .B(G832GAT_321_gat), .Y(G899GAT_329_gat) );
AND2XL U_g290 (.A(G831GAT_314_gat), .B(G830GAT_322_gat), .Y(G912GAT_330_gat) );
AND2XL U_g291 (.A(G829GAT_315_gat), .B(G828GAT_323_gat), .Y(G886GAT_331_gat) );
AND2XL U_g292 (.A(G827GAT_316_gat), .B(G826GAT_324_gat), .Y(G925GAT_332_gat) );
AND2XL U_g293 (.A(G825GAT_317_gat), .B(G824GAT_325_gat), .Y(G873GAT_333_gat) );
AND2XL U_g294 (.A(G823GAT_318_gat), .B(G822GAT_326_gat), .Y(G860GAT_334_gat) );
AND2XL U_g295 (.A(G821GAT_319_gat), .B(G820GAT_327_gat), .Y(G847GAT_335_gat) );
AND2XL U_g296 (.A(G819GAT_320_gat), .B(G818GAT_328_gat), .Y(G834GAT_336_gat) );
BUFX20 U_g297 (.A(G899GAT_329_gat), .Y(G951GAT_337_gat) );
BUFX20 U_g298 (.A(G899GAT_329_gat), .Y(G955GAT_338_gat) );
BUFX20 U_g299 (.A(G899GAT_329_gat), .Y(G963GAT_339_gat) );
BUFX20 U_g300 (.A(G899GAT_329_gat), .Y(G966GAT_340_gat) );
BUFX20 U_g301 (.A(G899GAT_329_gat), .Y(G969GAT_341_gat) );
BUFX20 U_g302 (.A(G912GAT_330_gat), .Y(G953GAT_342_gat) );
BUFX20 U_g303 (.A(G912GAT_330_gat), .Y(G957GAT_343_gat) );
BUFX20 U_g304 (.A(G912GAT_330_gat), .Y(G960GAT_344_gat) );
BUFX20 U_g305 (.A(G912GAT_330_gat), .Y(G965GAT_345_gat) );
BUFX20 U_g306 (.A(G912GAT_330_gat), .Y(G968GAT_346_gat) );
BUFX20 U_g307 (.A(G886GAT_331_gat), .Y(G950GAT_347_gat) );
BUFX20 U_g308 (.A(G886GAT_331_gat), .Y(G952GAT_348_gat) );
BUFX20 U_g309 (.A(G886GAT_331_gat), .Y(G959GAT_349_gat) );
BUFX20 U_g310 (.A(G886GAT_331_gat), .Y(G962GAT_350_gat) );
BUFX20 U_g311 (.A(G886GAT_331_gat), .Y(G967GAT_351_gat) );
BUFX20 U_g312 (.A(G925GAT_332_gat), .Y(G954GAT_352_gat) );
BUFX20 U_g313 (.A(G925GAT_332_gat), .Y(G956GAT_353_gat) );
BUFX20 U_g314 (.A(G925GAT_332_gat), .Y(G958GAT_354_gat) );
BUFX20 U_g315 (.A(G925GAT_332_gat), .Y(G961GAT_355_gat) );
BUFX20 U_g316 (.A(G925GAT_332_gat), .Y(G964GAT_356_gat) );
BUFX20 U_g317 (.A(G873GAT_333_gat), .Y(G943GAT_357_gat) );
BUFX20 U_g318 (.A(G873GAT_333_gat), .Y(G946GAT_358_gat) );
BUFX20 U_g319 (.A(G873GAT_333_gat), .Y(G949GAT_359_gat) );
BUFX20 U_g320 (.A(G873GAT_333_gat), .Y(G971GAT_360_gat) );
BUFX20 U_g321 (.A(G873GAT_333_gat), .Y(G975GAT_361_gat) );
BUFX20 U_g322 (.A(G860GAT_334_gat), .Y(G940GAT_362_gat) );
BUFX20 U_g323 (.A(G860GAT_334_gat), .Y(G945GAT_363_gat) );
BUFX20 U_g324 (.A(G860GAT_334_gat), .Y(G948GAT_364_gat) );
BUFX20 U_g325 (.A(G860GAT_334_gat), .Y(G973GAT_365_gat) );
BUFX20 U_g326 (.A(G860GAT_334_gat), .Y(G977GAT_366_gat) );
BUFX20 U_g327 (.A(G847GAT_335_gat), .Y(G939GAT_367_gat) );
BUFX20 U_g328 (.A(G847GAT_335_gat), .Y(G942GAT_368_gat) );
BUFX20 U_g329 (.A(G847GAT_335_gat), .Y(G947GAT_369_gat) );
BUFX20 U_g330 (.A(G847GAT_335_gat), .Y(G970GAT_370_gat) );
BUFX20 U_g331 (.A(G847GAT_335_gat), .Y(G972GAT_371_gat) );
BUFX20 U_g332 (.A(G834GAT_336_gat), .Y(G938GAT_372_gat) );
BUFX20 U_g333 (.A(G834GAT_336_gat), .Y(G941GAT_373_gat) );
BUFX20 U_g334 (.A(G834GAT_336_gat), .Y(G944GAT_374_gat) );
BUFX20 U_g335 (.A(G834GAT_336_gat), .Y(G974GAT_375_gat) );
BUFX20 U_g336 (.A(G834GAT_336_gat), .Y(G976GAT_376_gat) );
AND4XL U_g337 (.A(G899GAT_329_gat), .B(G960GAT_344_gat), .C(G959GAT_349_gat), .D(G958GAT_354_gat), .Y(G982GAT_377_gat) );
AND4XL U_g338 (.A(G963GAT_339_gat), .B(G912GAT_330_gat), .C(G962GAT_350_gat), .D(G961GAT_355_gat), .Y(G983GAT_378_gat) );
AND4XL U_g339 (.A(G966GAT_340_gat), .B(G965GAT_345_gat), .C(G886GAT_331_gat), .D(G964GAT_356_gat), .Y(G984GAT_379_gat) );
AND4XL U_g340 (.A(G969GAT_341_gat), .B(G968GAT_346_gat), .C(G967GAT_351_gat), .D(G925GAT_332_gat), .Y(G985GAT_380_gat) );
AND4XL U_g341 (.A(G873GAT_333_gat), .B(G940GAT_362_gat), .C(G939GAT_367_gat), .D(G938GAT_372_gat), .Y(G978GAT_381_gat) );
AND4XL U_g342 (.A(G943GAT_357_gat), .B(G860GAT_334_gat), .C(G942GAT_368_gat), .D(G941GAT_373_gat), .Y(G979GAT_382_gat) );
AND4XL U_g343 (.A(G946GAT_358_gat), .B(G945GAT_363_gat), .C(G847GAT_335_gat), .D(G944GAT_374_gat), .Y(G980GAT_383_gat) );
AND4XL U_g344 (.A(G949GAT_359_gat), .B(G948GAT_364_gat), .C(G947GAT_369_gat), .D(G834GAT_336_gat), .Y(G981GAT_384_gat) );
AND4XL U_g345 (.A(G985GAT_380_ngat), .B(G984GAT_379_ngat), .C(G983GAT_378_ngat), .D(G982GAT_377_ngat), .Y(G991GAT_385_gat) );
AND4XL U_g346 (.A(G981GAT_384_ngat), .B(G980GAT_383_ngat), .C(G979GAT_382_ngat), .D(G978GAT_381_ngat), .Y(G986GAT_386_gat) );
AND5XL U_g347 (.A(G986GAT_386_gat), .B(G899GAT_329_gat), .C(G953GAT_342_gat), .D(G952GAT_348_gat), .E(G925GAT_332_gat), .Y(G1001GAT_387_gat) );
AND5XL U_g348 (.A(G986GAT_386_gat), .B(G899GAT_329_gat), .C(G957GAT_343_gat), .D(G886GAT_331_gat), .E(G956GAT_353_gat), .Y(G1011GAT_388_gat) );
AND5XL U_g349 (.A(G986GAT_386_gat), .B(G951GAT_337_gat), .C(G912GAT_330_gat), .D(G950GAT_347_gat), .E(G925GAT_332_gat), .Y(G996GAT_389_gat) );
AND5XL U_g350 (.A(G986GAT_386_gat), .B(G955GAT_338_gat), .C(G912GAT_330_gat), .D(G886GAT_331_gat), .E(G954GAT_352_gat), .Y(G1006GAT_390_gat) );
AND5XL U_g351 (.A(G991GAT_385_gat), .B(G873GAT_333_gat), .C(G973GAT_365_gat), .D(G972GAT_371_gat), .E(G834GAT_336_gat), .Y(G1021GAT_391_gat) );
AND5XL U_g352 (.A(G991GAT_385_gat), .B(G873GAT_333_gat), .C(G977GAT_366_gat), .D(G847GAT_335_gat), .E(G976GAT_376_gat), .Y(G1031GAT_392_gat) );
AND5XL U_g353 (.A(G991GAT_385_gat), .B(G971GAT_360_gat), .C(G860GAT_334_gat), .D(G970GAT_370_gat), .E(G834GAT_336_gat), .Y(G1016GAT_393_gat) );
AND5XL U_g354 (.A(G991GAT_385_gat), .B(G975GAT_361_gat), .C(G860GAT_334_gat), .D(G847GAT_335_gat), .E(G974GAT_375_gat), .Y(G1026GAT_394_gat) );
AND2XL U_g355 (.A(G1016GAT_393_gat), .B(G899GAT_329_gat), .Y(G1093GAT_395_gat) );
AND2XL U_g356 (.A(G1021GAT_391_gat), .B(G899GAT_329_gat), .Y(G1105GAT_396_gat) );
AND2XL U_g357 (.A(G1026GAT_394_gat), .B(G899GAT_329_gat), .Y(G1117GAT_397_gat) );
AND2XL U_g358 (.A(G1031GAT_392_gat), .B(G899GAT_329_gat), .Y(G1129GAT_398_gat) );
AND2XL U_g359 (.A(G1016GAT_393_gat), .B(G912GAT_330_gat), .Y(G1090GAT_399_gat) );
AND2XL U_g360 (.A(G1021GAT_391_gat), .B(G912GAT_330_gat), .Y(G1102GAT_400_gat) );
AND2XL U_g361 (.A(G1026GAT_394_gat), .B(G912GAT_330_gat), .Y(G1114GAT_401_gat) );
AND2XL U_g362 (.A(G1031GAT_392_gat), .B(G912GAT_330_gat), .Y(G1126GAT_402_gat) );
AND2XL U_g363 (.A(G1016GAT_393_gat), .B(G886GAT_331_gat), .Y(G1087GAT_403_gat) );
AND2XL U_g364 (.A(G1021GAT_391_gat), .B(G886GAT_331_gat), .Y(G1099GAT_404_gat) );
AND2XL U_g365 (.A(G1026GAT_394_gat), .B(G886GAT_331_gat), .Y(G1111GAT_405_gat) );
AND2XL U_g366 (.A(G1031GAT_392_gat), .B(G886GAT_331_gat), .Y(G1123GAT_406_gat) );
AND2XL U_g367 (.A(G1016GAT_393_gat), .B(G925GAT_332_gat), .Y(G1084GAT_407_gat) );
AND2XL U_g368 (.A(G1021GAT_391_gat), .B(G925GAT_332_gat), .Y(G1096GAT_408_gat) );
AND2XL U_g369 (.A(G1026GAT_394_gat), .B(G925GAT_332_gat), .Y(G1108GAT_409_gat) );
AND2XL U_g370 (.A(G1031GAT_392_gat), .B(G925GAT_332_gat), .Y(G1120GAT_410_gat) );
AND2XL U_g371 (.A(G996GAT_389_gat), .B(G873GAT_333_gat), .Y(G1045GAT_411_gat) );
AND2XL U_g372 (.A(G1001GAT_387_gat), .B(G873GAT_333_gat), .Y(G1057GAT_412_gat) );
AND2XL U_g373 (.A(G1006GAT_390_gat), .B(G873GAT_333_gat), .Y(G1069GAT_413_gat) );
AND2XL U_g374 (.A(G1011GAT_388_gat), .B(G873GAT_333_gat), .Y(G1081GAT_414_gat) );
AND2XL U_g375 (.A(G996GAT_389_gat), .B(G860GAT_334_gat), .Y(G1042GAT_415_gat) );
AND2XL U_g376 (.A(G1001GAT_387_gat), .B(G860GAT_334_gat), .Y(G1054GAT_416_gat) );
AND2XL U_g377 (.A(G1006GAT_390_gat), .B(G860GAT_334_gat), .Y(G1066GAT_417_gat) );
AND2XL U_g378 (.A(G1011GAT_388_gat), .B(G860GAT_334_gat), .Y(G1078GAT_418_gat) );
AND2XL U_g379 (.A(G996GAT_389_gat), .B(G847GAT_335_gat), .Y(G1039GAT_419_gat) );
AND2XL U_g380 (.A(G1001GAT_387_gat), .B(G847GAT_335_gat), .Y(G1051GAT_420_gat) );
AND2XL U_g381 (.A(G1006GAT_390_gat), .B(G847GAT_335_gat), .Y(G1063GAT_421_gat) );
AND2XL U_g382 (.A(G1011GAT_388_gat), .B(G847GAT_335_gat), .Y(G1075GAT_422_gat) );
AND2XL U_g383 (.A(G996GAT_389_gat), .B(G834GAT_336_gat), .Y(G1036GAT_423_gat) );
AND2XL U_g384 (.A(G1001GAT_387_gat), .B(G834GAT_336_gat), .Y(G1048GAT_424_gat) );
AND2XL U_g385 (.A(G1006GAT_390_gat), .B(G834GAT_336_gat), .Y(G1060GAT_425_gat) );
AND2XL U_g386 (.A(G1011GAT_388_gat), .B(G834GAT_336_gat), .Y(G1072GAT_426_gat) );
AND2XL U_g387 (.A(G1129GAT_398_gat), .B(G218GAT_31_gat), .Y(G1225GAT_427_gat) );
AND2XL U_g388 (.A(G1126GAT_402_gat), .B(G211GAT_30_gat), .Y(G1222GAT_428_gat) );
AND2XL U_g389 (.A(G1123GAT_406_gat), .B(G204GAT_29_gat), .Y(G1219GAT_429_gat) );
AND2XL U_g390 (.A(G1120GAT_410_gat), .B(G197GAT_28_gat), .Y(G1216GAT_430_gat) );
AND2XL U_g391 (.A(G1117GAT_397_gat), .B(G190GAT_27_gat), .Y(G1213GAT_431_gat) );
AND2XL U_g392 (.A(G1114GAT_401_gat), .B(G183GAT_26_gat), .Y(G1210GAT_432_gat) );
AND2XL U_g393 (.A(G1111GAT_405_gat), .B(G176GAT_25_gat), .Y(G1207GAT_433_gat) );
AND2XL U_g394 (.A(G1108GAT_409_gat), .B(G169GAT_24_gat), .Y(G1204GAT_434_gat) );
AND2XL U_g395 (.A(G1105GAT_396_gat), .B(G162GAT_23_gat), .Y(G1201GAT_435_gat) );
AND2XL U_g396 (.A(G1102GAT_400_gat), .B(G155GAT_22_gat), .Y(G1198GAT_436_gat) );
AND2XL U_g397 (.A(G1099GAT_404_gat), .B(G148GAT_21_gat), .Y(G1195GAT_437_gat) );
AND2XL U_g398 (.A(G1096GAT_408_gat), .B(G141GAT_20_gat), .Y(G1192GAT_438_gat) );
AND2XL U_g399 (.A(G1093GAT_395_gat), .B(G134GAT_19_gat), .Y(G1189GAT_439_gat) );
AND2XL U_g400 (.A(G1090GAT_399_gat), .B(G127GAT_18_gat), .Y(G1186GAT_440_gat) );
AND2XL U_g401 (.A(G1087GAT_403_gat), .B(G120GAT_17_gat), .Y(G1183GAT_441_gat) );
AND2XL U_g402 (.A(G1084GAT_407_gat), .B(G113GAT_16_gat), .Y(G1180GAT_442_gat) );
AND2XL U_g403 (.A(G1081GAT_414_gat), .B(G106GAT_15_gat), .Y(G1177GAT_443_gat) );
AND2XL U_g404 (.A(G1078GAT_418_gat), .B(G99GAT_14_gat), .Y(G1174GAT_444_gat) );
AND2XL U_g405 (.A(G1075GAT_422_gat), .B(G92GAT_13_gat), .Y(G1171GAT_445_gat) );
AND2XL U_g406 (.A(G1072GAT_426_gat), .B(G85GAT_12_gat), .Y(G1168GAT_446_gat) );
AND2XL U_g407 (.A(G1069GAT_413_gat), .B(G78GAT_11_gat), .Y(G1165GAT_447_gat) );
AND2XL U_g408 (.A(G1066GAT_417_gat), .B(G71GAT_10_gat), .Y(G1162GAT_448_gat) );
AND2XL U_g409 (.A(G1063GAT_421_gat), .B(G64GAT_9_gat), .Y(G1159GAT_449_gat) );
AND2XL U_g410 (.A(G1060GAT_425_gat), .B(G57GAT_8_gat), .Y(G1156GAT_450_gat) );
AND2XL U_g411 (.A(G1057GAT_412_gat), .B(G50GAT_7_gat), .Y(G1153GAT_451_gat) );
AND2XL U_g412 (.A(G1054GAT_416_gat), .B(G43GAT_6_gat), .Y(G1150GAT_452_gat) );
AND2XL U_g413 (.A(G1051GAT_420_gat), .B(G36GAT_5_gat), .Y(G1147GAT_453_gat) );
AND2XL U_g414 (.A(G1048GAT_424_gat), .B(G29GAT_4_gat), .Y(G1144GAT_454_gat) );
AND2XL U_g415 (.A(G1045GAT_411_gat), .B(G22GAT_3_gat), .Y(G1141GAT_455_gat) );
AND2XL U_g416 (.A(G1042GAT_415_gat), .B(G15GAT_2_gat), .Y(G1138GAT_456_gat) );
AND2XL U_g417 (.A(G1039GAT_419_gat), .B(G8GAT_1_gat), .Y(G1135GAT_457_gat) );
AND2XL U_g418 (.A(G1036GAT_423_gat), .B(G1GAT_0_gat), .Y(G1132GAT_458_gat) );
AND2XL U_g419 (.A(G1189GAT_439_gat), .B(G1093GAT_395_gat), .Y(G1267GAT_459_gat) );
AND2XL U_g420 (.A(G1201GAT_435_gat), .B(G1105GAT_396_gat), .Y(G1275GAT_460_gat) );
AND2XL U_g421 (.A(G1213GAT_431_gat), .B(G1117GAT_397_gat), .Y(G1283GAT_461_gat) );
AND2XL U_g422 (.A(G1225GAT_427_gat), .B(G1129GAT_398_gat), .Y(G1291GAT_462_gat) );
AND2XL U_g423 (.A(G1186GAT_440_gat), .B(G1090GAT_399_gat), .Y(G1265GAT_463_gat) );
AND2XL U_g424 (.A(G1198GAT_436_gat), .B(G1102GAT_400_gat), .Y(G1273GAT_464_gat) );
AND2XL U_g425 (.A(G1210GAT_432_gat), .B(G1114GAT_401_gat), .Y(G1281GAT_465_gat) );
AND2XL U_g426 (.A(G1222GAT_428_gat), .B(G1126GAT_402_gat), .Y(G1289GAT_466_gat) );
AND2XL U_g427 (.A(G1183GAT_441_gat), .B(G1087GAT_403_gat), .Y(G1263GAT_467_gat) );
AND2XL U_g428 (.A(G1195GAT_437_gat), .B(G1099GAT_404_gat), .Y(G1271GAT_468_gat) );
AND2XL U_g429 (.A(G1207GAT_433_gat), .B(G1111GAT_405_gat), .Y(G1279GAT_469_gat) );
AND2XL U_g430 (.A(G1219GAT_429_gat), .B(G1123GAT_406_gat), .Y(G1287GAT_470_gat) );
AND2XL U_g431 (.A(G1180GAT_442_gat), .B(G1084GAT_407_gat), .Y(G1261GAT_471_gat) );
AND2XL U_g432 (.A(G1192GAT_438_gat), .B(G1096GAT_408_gat), .Y(G1269GAT_472_gat) );
AND2XL U_g433 (.A(G1204GAT_434_gat), .B(G1108GAT_409_gat), .Y(G1277GAT_473_gat) );
AND2XL U_g434 (.A(G1216GAT_430_gat), .B(G1120GAT_410_gat), .Y(G1285GAT_474_gat) );
AND2XL U_g435 (.A(G1141GAT_455_gat), .B(G1045GAT_411_gat), .Y(G1235GAT_475_gat) );
AND2XL U_g436 (.A(G1153GAT_451_gat), .B(G1057GAT_412_gat), .Y(G1243GAT_476_gat) );
AND2XL U_g437 (.A(G1165GAT_447_gat), .B(G1069GAT_413_gat), .Y(G1251GAT_477_gat) );
AND2XL U_g438 (.A(G1177GAT_443_gat), .B(G1081GAT_414_gat), .Y(G1259GAT_478_gat) );
AND2XL U_g439 (.A(G1138GAT_456_gat), .B(G1042GAT_415_gat), .Y(G1233GAT_479_gat) );
AND2XL U_g440 (.A(G1150GAT_452_gat), .B(G1054GAT_416_gat), .Y(G1241GAT_480_gat) );
AND2XL U_g441 (.A(G1162GAT_448_gat), .B(G1066GAT_417_gat), .Y(G1249GAT_481_gat) );
AND2XL U_g442 (.A(G1174GAT_444_gat), .B(G1078GAT_418_gat), .Y(G1257GAT_482_gat) );
AND2XL U_g443 (.A(G1135GAT_457_gat), .B(G1039GAT_419_gat), .Y(G1231GAT_483_gat) );
AND2XL U_g444 (.A(G1147GAT_453_gat), .B(G1051GAT_420_gat), .Y(G1239GAT_484_gat) );
AND2XL U_g445 (.A(G1159GAT_449_gat), .B(G1063GAT_421_gat), .Y(G1247GAT_485_gat) );
AND2XL U_g446 (.A(G1171GAT_445_gat), .B(G1075GAT_422_gat), .Y(G1255GAT_486_gat) );
AND2XL U_g447 (.A(G1132GAT_458_gat), .B(G1036GAT_423_gat), .Y(G1229GAT_487_gat) );
AND2XL U_g448 (.A(G1144GAT_454_gat), .B(G1048GAT_424_gat), .Y(G1237GAT_488_gat) );
AND2XL U_g449 (.A(G1156GAT_450_gat), .B(G1060GAT_425_gat), .Y(G1245GAT_489_gat) );
AND2XL U_g450 (.A(G1168GAT_446_gat), .B(G1072GAT_426_gat), .Y(G1253GAT_490_gat) );
AND2XL U_g451 (.A(G1225GAT_427_gat), .B(G218GAT_31_gat), .Y(G1290GAT_491_gat) );
AND2XL U_g452 (.A(G1222GAT_428_gat), .B(G211GAT_30_gat), .Y(G1288GAT_492_gat) );
AND2XL U_g453 (.A(G1219GAT_429_gat), .B(G204GAT_29_gat), .Y(G1286GAT_493_gat) );
AND2XL U_g454 (.A(G1216GAT_430_gat), .B(G197GAT_28_gat), .Y(G1284GAT_494_gat) );
AND2XL U_g455 (.A(G1213GAT_431_gat), .B(G190GAT_27_gat), .Y(G1282GAT_495_gat) );
AND2XL U_g456 (.A(G1210GAT_432_gat), .B(G183GAT_26_gat), .Y(G1280GAT_496_gat) );
AND2XL U_g457 (.A(G1207GAT_433_gat), .B(G176GAT_25_gat), .Y(G1278GAT_497_gat) );
AND2XL U_g458 (.A(G1204GAT_434_gat), .B(G169GAT_24_gat), .Y(G1276GAT_498_gat) );
AND2XL U_g459 (.A(G1201GAT_435_gat), .B(G162GAT_23_gat), .Y(G1274GAT_499_gat) );
AND2XL U_g460 (.A(G1198GAT_436_gat), .B(G155GAT_22_gat), .Y(G1272GAT_500_gat) );
AND2XL U_g461 (.A(G1195GAT_437_gat), .B(G148GAT_21_gat), .Y(G1270GAT_501_gat) );
AND2XL U_g462 (.A(G1192GAT_438_gat), .B(G141GAT_20_gat), .Y(G1268GAT_502_gat) );
AND2XL U_g463 (.A(G1189GAT_439_gat), .B(G134GAT_19_gat), .Y(G1266GAT_503_gat) );
AND2XL U_g464 (.A(G1186GAT_440_gat), .B(G127GAT_18_gat), .Y(G1264GAT_504_gat) );
AND2XL U_g465 (.A(G1183GAT_441_gat), .B(G120GAT_17_gat), .Y(G1262GAT_505_gat) );
AND2XL U_g466 (.A(G1180GAT_442_gat), .B(G113GAT_16_gat), .Y(G1260GAT_506_gat) );
AND2XL U_g467 (.A(G1177GAT_443_gat), .B(G106GAT_15_gat), .Y(G1258GAT_507_gat) );
AND2XL U_g468 (.A(G1174GAT_444_gat), .B(G99GAT_14_gat), .Y(G1256GAT_508_gat) );
AND2XL U_g469 (.A(G1171GAT_445_gat), .B(G92GAT_13_gat), .Y(G1254GAT_509_gat) );
AND2XL U_g470 (.A(G1168GAT_446_gat), .B(G85GAT_12_gat), .Y(G1252GAT_510_gat) );
AND2XL U_g471 (.A(G1165GAT_447_gat), .B(G78GAT_11_gat), .Y(G1250GAT_511_gat) );
AND2XL U_g472 (.A(G1162GAT_448_gat), .B(G71GAT_10_gat), .Y(G1248GAT_512_gat) );
AND2XL U_g473 (.A(G1159GAT_449_gat), .B(G64GAT_9_gat), .Y(G1246GAT_513_gat) );
AND2XL U_g474 (.A(G1156GAT_450_gat), .B(G57GAT_8_gat), .Y(G1244GAT_514_gat) );
AND2XL U_g475 (.A(G1153GAT_451_gat), .B(G50GAT_7_gat), .Y(G1242GAT_515_gat) );
AND2XL U_g476 (.A(G1150GAT_452_gat), .B(G43GAT_6_gat), .Y(G1240GAT_516_gat) );
AND2XL U_g477 (.A(G1147GAT_453_gat), .B(G36GAT_5_gat), .Y(G1238GAT_517_gat) );
AND2XL U_g478 (.A(G1144GAT_454_gat), .B(G29GAT_4_gat), .Y(G1236GAT_518_gat) );
AND2XL U_g479 (.A(G1141GAT_455_gat), .B(G22GAT_3_gat), .Y(G1234GAT_519_gat) );
AND2XL U_g480 (.A(G1138GAT_456_gat), .B(G15GAT_2_gat), .Y(G1232GAT_520_gat) );
AND2XL U_g481 (.A(G1135GAT_457_gat), .B(G8GAT_1_gat), .Y(G1230GAT_521_gat) );
AND2XL U_g482 (.A(G1132GAT_458_gat), .B(G1GAT_0_gat), .Y(G1228GAT_522_gat) );
AND2XL U_g483 (.A(G1267GAT_459_gat), .B(G1266GAT_503_gat), .Y(G1311GAT_523_gat) );
AND2XL U_g484 (.A(G1275GAT_460_gat), .B(G1274GAT_499_gat), .Y(G1315GAT_524_gat) );
AND2XL U_g485 (.A(G1283GAT_461_gat), .B(G1282GAT_495_gat), .Y(G1319GAT_525_gat) );
AND2XL U_g486 (.A(G1291GAT_462_gat), .B(G1290GAT_491_gat), .Y(G1323GAT_526_gat) );
AND2XL U_g487 (.A(G1265GAT_463_gat), .B(G1264GAT_504_gat), .Y(G1310GAT_527_gat) );
AND2XL U_g488 (.A(G1273GAT_464_gat), .B(G1272GAT_500_gat), .Y(G1314GAT_528_gat) );
AND2XL U_g489 (.A(G1281GAT_465_gat), .B(G1280GAT_496_gat), .Y(G1318GAT_529_gat) );
AND2XL U_g490 (.A(G1289GAT_466_gat), .B(G1288GAT_492_gat), .Y(G1322GAT_530_gat) );
AND2XL U_g491 (.A(G1263GAT_467_gat), .B(G1262GAT_505_gat), .Y(G1309GAT_531_gat) );
AND2XL U_g492 (.A(G1271GAT_468_gat), .B(G1270GAT_501_gat), .Y(G1313GAT_532_gat) );
AND2XL U_g493 (.A(G1279GAT_469_gat), .B(G1278GAT_497_gat), .Y(G1317GAT_533_gat) );
AND2XL U_g494 (.A(G1287GAT_470_gat), .B(G1286GAT_493_gat), .Y(G1321GAT_534_gat) );
AND2XL U_g495 (.A(G1261GAT_471_gat), .B(G1260GAT_506_gat), .Y(G1308GAT_535_gat) );
AND2XL U_g496 (.A(G1269GAT_472_gat), .B(G1268GAT_502_gat), .Y(G1312GAT_536_gat) );
AND2XL U_g497 (.A(G1277GAT_473_gat), .B(G1276GAT_498_gat), .Y(G1316GAT_537_gat) );
AND2XL U_g498 (.A(G1285GAT_474_gat), .B(G1284GAT_494_gat), .Y(G1320GAT_538_gat) );
AND2XL U_g499 (.A(G1235GAT_475_gat), .B(G1234GAT_519_gat), .Y(G1295GAT_539_gat) );
AND2XL U_g500 (.A(G1243GAT_476_gat), .B(G1242GAT_515_gat), .Y(G1299GAT_540_gat) );
AND2XL U_g501 (.A(G1251GAT_477_gat), .B(G1250GAT_511_gat), .Y(G1303GAT_541_gat) );
AND2XL U_g502 (.A(G1259GAT_478_gat), .B(G1258GAT_507_gat), .Y(G1307GAT_542_gat) );
AND2XL U_g503 (.A(G1233GAT_479_gat), .B(G1232GAT_520_gat), .Y(G1294GAT_543_gat) );
AND2XL U_g504 (.A(G1241GAT_480_gat), .B(G1240GAT_516_gat), .Y(G1298GAT_544_gat) );
AND2XL U_g505 (.A(G1249GAT_481_gat), .B(G1248GAT_512_gat), .Y(G1302GAT_545_gat) );
AND2XL U_g506 (.A(G1257GAT_482_gat), .B(G1256GAT_508_gat), .Y(G1306GAT_546_gat) );
AND2XL U_g507 (.A(G1231GAT_483_gat), .B(G1230GAT_521_gat), .Y(G1293GAT_547_gat) );
AND2XL U_g508 (.A(G1239GAT_484_gat), .B(G1238GAT_517_gat), .Y(G1297GAT_548_gat) );
AND2XL U_g509 (.A(G1247GAT_485_gat), .B(G1246GAT_513_gat), .Y(G1301GAT_549_gat) );
AND2XL U_g510 (.A(G1255GAT_486_gat), .B(G1254GAT_509_gat), .Y(G1305GAT_550_gat) );
AND2XL U_g511 (.A(G1229GAT_487_gat), .B(G1228GAT_522_gat), .Y(G1292GAT_551_gat) );
AND2XL U_g512 (.A(G1237GAT_488_gat), .B(G1236GAT_518_gat), .Y(G1296GAT_552_gat) );
AND2XL U_g513 (.A(G1245GAT_489_gat), .B(G1244GAT_514_gat), .Y(G1300GAT_553_gat) );
AND2XL U_g514 (.A(G1253GAT_490_gat), .B(G1252GAT_510_gat), .Y(G1304GAT_554_gat) );
BUFX20 U_g515 (.A(G1311GAT_523_gat), .Y(G1343GAT_555_gat) );
BUFX20 U_g516 (.A(G1315GAT_524_gat), .Y(G1347GAT_556_gat) );
BUFX20 U_g517 (.A(G1319GAT_525_gat), .Y(G1351GAT_557_gat) );
BUFX20 U_g518 (.A(G1323GAT_526_gat), .Y(G1355GAT_558_gat) );
BUFX20 U_g519 (.A(G1310GAT_527_gat), .Y(G1342GAT_559_gat) );
BUFX20 U_g520 (.A(G1314GAT_528_gat), .Y(G1346GAT_560_gat) );
BUFX20 U_g521 (.A(G1318GAT_529_gat), .Y(G1350GAT_561_gat) );
BUFX20 U_g522 (.A(G1322GAT_530_gat), .Y(G1354GAT_562_gat) );
BUFX20 U_g523 (.A(G1309GAT_531_gat), .Y(G1341GAT_563_gat) );
BUFX20 U_g524 (.A(G1313GAT_532_gat), .Y(G1345GAT_564_gat) );
BUFX20 U_g525 (.A(G1317GAT_533_gat), .Y(G1349GAT_565_gat) );
BUFX20 U_g526 (.A(G1321GAT_534_gat), .Y(G1353GAT_566_gat) );
BUFX20 U_g527 (.A(G1308GAT_535_gat), .Y(G1340GAT_567_gat) );
BUFX20 U_g528 (.A(G1312GAT_536_gat), .Y(G1344GAT_568_gat) );
BUFX20 U_g529 (.A(G1316GAT_537_gat), .Y(G1348GAT_569_gat) );
BUFX20 U_g530 (.A(G1320GAT_538_gat), .Y(G1352GAT_570_gat) );
BUFX20 U_g531 (.A(G1295GAT_539_gat), .Y(G1327GAT_571_gat) );
BUFX20 U_g532 (.A(G1299GAT_540_gat), .Y(G1331GAT_572_gat) );
BUFX20 U_g533 (.A(G1303GAT_541_gat), .Y(G1335GAT_573_gat) );
BUFX20 U_g534 (.A(G1307GAT_542_gat), .Y(G1339GAT_574_gat) );
BUFX20 U_g535 (.A(G1294GAT_543_gat), .Y(G1326GAT_575_gat) );
BUFX20 U_g536 (.A(G1298GAT_544_gat), .Y(G1330GAT_576_gat) );
BUFX20 U_g537 (.A(G1302GAT_545_gat), .Y(G1334GAT_577_gat) );
BUFX20 U_g538 (.A(G1306GAT_546_gat), .Y(G1338GAT_578_gat) );
BUFX20 U_g539 (.A(G1293GAT_547_gat), .Y(G1325GAT_579_gat) );
BUFX20 U_g540 (.A(G1297GAT_548_gat), .Y(G1329GAT_580_gat) );
BUFX20 U_g541 (.A(G1301GAT_549_gat), .Y(G1333GAT_581_gat) );
BUFX20 U_g542 (.A(G1305GAT_550_gat), .Y(G1337GAT_582_gat) );
BUFX20 U_g543 (.A(G1292GAT_551_gat), .Y(G1324GAT_583_gat) );
BUFX20 U_g544 (.A(G1296GAT_552_gat), .Y(G1328GAT_584_gat) );
BUFX20 U_g545 (.A(G1300GAT_553_gat), .Y(G1332GAT_585_gat) );
BUFX20 U_g546 (.A(G1304GAT_554_gat), .Y(G1336GAT_586_gat) );
INVXL U_g547 (.A(G982GAT_377_gat), .Y(G982GAT_377_ngat) );
INVXL U_g548 (.A(G983GAT_378_gat), .Y(G983GAT_378_ngat) );
INVXL U_g549 (.A(G984GAT_379_gat), .Y(G984GAT_379_ngat) );
INVXL U_g550 (.A(G985GAT_380_gat), .Y(G985GAT_380_ngat) );
INVXL U_g551 (.A(G978GAT_381_gat), .Y(G978GAT_381_ngat) );
INVXL U_g552 (.A(G979GAT_382_gat), .Y(G979GAT_382_ngat) );
INVXL U_g553 (.A(G980GAT_383_gat), .Y(G980GAT_383_ngat) );
INVXL U_g554 (.A(G981GAT_384_gat), .Y(G981GAT_384_ngat) );

endmodule
