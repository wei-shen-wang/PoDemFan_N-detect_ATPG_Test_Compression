module C432 ( G1GAT_0_gat, G4GAT_1_gat, G8GAT_2_gat, G11GAT_3_gat, G14GAT_4_gat, G17GAT_5_gat, G21GAT_6_gat, G24GAT_7_gat, G27GAT_8_gat, G30GAT_9_gat, G34GAT_10_gat, G37GAT_11_gat, G40GAT_12_gat, G43GAT_13_gat, G47GAT_14_gat, G50GAT_15_gat, G53GAT_16_gat, G56GAT_17_gat, G60GAT_18_gat, G63GAT_19_gat, G66GAT_20_gat, G69GAT_21_gat, G73GAT_22_gat, G76GAT_23_gat, G79GAT_24_gat, G82GAT_25_gat, G86GAT_26_gat, G89GAT_27_gat, G92GAT_28_gat, G95GAT_29_gat, G99GAT_30_gat, G102GAT_31_gat, G105GAT_32_gat, G108GAT_33_gat, G112GAT_34_gat, G115GAT_35_gat, G223GAT_84_gat, G329GAT_133_gat, G370GAT_163_gat, G421GAT_188_gat, G430GAT_193_gat, G431GAT_194_gat, G432GAT_195_gat);

input G1GAT_0_gat;
input G4GAT_1_gat;
input G8GAT_2_gat;
input G11GAT_3_gat;
input G14GAT_4_gat;
input G17GAT_5_gat;
input G21GAT_6_gat;
input G24GAT_7_gat;
input G27GAT_8_gat;
input G30GAT_9_gat;
input G34GAT_10_gat;
input G37GAT_11_gat;
input G40GAT_12_gat;
input G43GAT_13_gat;
input G47GAT_14_gat;
input G50GAT_15_gat;
input G53GAT_16_gat;
input G56GAT_17_gat;
input G60GAT_18_gat;
input G63GAT_19_gat;
input G66GAT_20_gat;
input G69GAT_21_gat;
input G73GAT_22_gat;
input G76GAT_23_gat;
input G79GAT_24_gat;
input G82GAT_25_gat;
input G86GAT_26_gat;
input G89GAT_27_gat;
input G92GAT_28_gat;
input G95GAT_29_gat;
input G99GAT_30_gat;
input G102GAT_31_gat;
input G105GAT_32_gat;
input G108GAT_33_gat;
input G112GAT_34_gat;
input G115GAT_35_gat;

output G223GAT_84_gat;
output G329GAT_133_gat;
output G370GAT_163_gat;
output G421GAT_188_gat;
output G430GAT_193_gat;
output G431GAT_194_gat;
output G432GAT_195_gat;

BUFX20 U_g1 (.A(G108GAT_33_gat), .Y(G151GAT_36_gat) );
BUFX20 U_g2 (.A(G102GAT_31_gat), .Y(G150GAT_37_gat) );
BUFX20 U_g3 (.A(G95GAT_29_gat), .Y(G147GAT_38_gat) );
BUFX20 U_g4 (.A(G89GAT_27_gat), .Y(G146GAT_39_gat) );
BUFX20 U_g5 (.A(G82GAT_25_gat), .Y(G143GAT_40_gat) );
BUFX20 U_g6 (.A(G76GAT_23_gat), .Y(G142GAT_41_gat) );
BUFX20 U_g7 (.A(G69GAT_21_gat), .Y(G139GAT_42_gat) );
BUFX20 U_g8 (.A(G63GAT_19_gat), .Y(G138GAT_43_gat) );
BUFX20 U_g9 (.A(G56GAT_17_gat), .Y(G135GAT_44_gat) );
BUFX20 U_g10 (.A(G50GAT_15_gat), .Y(G134GAT_45_gat) );
BUFX20 U_g11 (.A(G43GAT_13_gat), .Y(G131GAT_46_gat) );
BUFX20 U_g12 (.A(G37GAT_11_gat), .Y(G130GAT_47_gat) );
BUFX20 U_g13 (.A(G30GAT_9_gat), .Y(G127GAT_48_gat) );
BUFX20 U_g14 (.A(G24GAT_7_gat), .Y(G126GAT_49_gat) );
BUFX20 U_g15 (.A(G17GAT_5_gat), .Y(G123GAT_50_gat) );
BUFX20 U_g16 (.A(G11GAT_3_gat), .Y(G122GAT_51_gat) );
BUFX20 U_g17 (.A(G4GAT_1_gat), .Y(G119GAT_52_gat) );
BUFX20 U_g18 (.A(G1GAT_0_gat), .Y(G118GAT_53_gat) );
AND2XL U_g19 (.A(G151GAT_36_ngat), .B(G115GAT_35_ngat), .Y(G198GAT_54_gat) );
AND2XL U_g20 (.A(G151GAT_36_ngat), .B(G112GAT_34_ngat), .Y(G197GAT_55_gat) );
AND2XL U_g21 (.A(G108GAT_33_gat), .B(G150GAT_37_gat), .Y(G180GAT_56_gat) );
AND2XL U_g22 (.A(G147GAT_38_ngat), .B(G105GAT_32_ngat), .Y(G196GAT_57_gat) );
AND2XL U_g23 (.A(G147GAT_38_ngat), .B(G99GAT_30_ngat), .Y(G195GAT_58_gat) );
AND2XL U_g24 (.A(G95GAT_29_gat), .B(G146GAT_39_gat), .Y(G177GAT_59_gat) );
AND2XL U_g25 (.A(G143GAT_40_ngat), .B(G92GAT_28_ngat), .Y(G194GAT_60_gat) );
AND2XL U_g26 (.A(G143GAT_40_ngat), .B(G86GAT_26_ngat), .Y(G193GAT_61_gat) );
AND2XL U_g27 (.A(G82GAT_25_gat), .B(G142GAT_41_gat), .Y(G174GAT_62_gat) );
AND2XL U_g28 (.A(G139GAT_42_ngat), .B(G79GAT_24_ngat), .Y(G192GAT_63_gat) );
AND2XL U_g29 (.A(G139GAT_42_ngat), .B(G73GAT_22_ngat), .Y(G191GAT_64_gat) );
AND2XL U_g30 (.A(G69GAT_21_gat), .B(G138GAT_43_gat), .Y(G171GAT_65_gat) );
AND2XL U_g31 (.A(G135GAT_44_ngat), .B(G66GAT_20_ngat), .Y(G190GAT_66_gat) );
AND2XL U_g32 (.A(G135GAT_44_ngat), .B(G60GAT_18_ngat), .Y(G189GAT_67_gat) );
AND2XL U_g33 (.A(G56GAT_17_gat), .B(G134GAT_45_gat), .Y(G168GAT_68_gat) );
AND2XL U_g34 (.A(G131GAT_46_ngat), .B(G53GAT_16_ngat), .Y(G188GAT_69_gat) );
AND2XL U_g35 (.A(G131GAT_46_ngat), .B(G47GAT_14_ngat), .Y(G187GAT_70_gat) );
AND2XL U_g36 (.A(G43GAT_13_gat), .B(G130GAT_47_gat), .Y(G165GAT_71_gat) );
AND2XL U_g37 (.A(G127GAT_48_ngat), .B(G40GAT_12_ngat), .Y(G186GAT_72_gat) );
AND2XL U_g38 (.A(G127GAT_48_ngat), .B(G34GAT_10_ngat), .Y(G185GAT_73_gat) );
AND2XL U_g39 (.A(G30GAT_9_gat), .B(G126GAT_49_gat), .Y(G162GAT_74_gat) );
AND2XL U_g40 (.A(G123GAT_50_ngat), .B(G27GAT_8_ngat), .Y(G184GAT_75_gat) );
AND2XL U_g41 (.A(G123GAT_50_ngat), .B(G21GAT_6_ngat), .Y(G183GAT_76_gat) );
AND2XL U_g42 (.A(G17GAT_5_gat), .B(G122GAT_51_gat), .Y(G159GAT_77_gat) );
AND2XL U_g43 (.A(G119GAT_52_ngat), .B(G14GAT_4_ngat), .Y(G158GAT_78_gat) );
AND2XL U_g44 (.A(G119GAT_52_ngat), .B(G8GAT_2_ngat), .Y(G157GAT_79_gat) );
AND2XL U_g45 (.A(G4GAT_1_gat), .B(G118GAT_53_gat), .Y(G154GAT_80_gat) );
AND9XL U_g46 (.A(G180GAT_56_gat), .B(G177GAT_59_gat), .C(G174GAT_62_gat), .D(G171GAT_65_gat), .E(G168GAT_68_gat), .F(G165GAT_71_gat), .G(G162GAT_74_gat), .H(G159GAT_77_gat), .I(G154GAT_80_gat), .Y(G199GAT_81_gat) );
BUFX20 U_g47 (.A(G199GAT_81_gat), .Y(G203GAT_82_gat) );
BUFX20 U_g48 (.A(G199GAT_81_gat), .Y(G213GAT_83_gat) );
BUFX20 U_g49 (.A(G199GAT_81_gat), .Y(G223GAT_84_gat) );
OR2XL U_g50 (.A(Ginternal__52gat), .B(Ginternal__51gat), .Y(G251GAT_85_gat) );
AND2XL U_g51 (.A(G180GAT_56_gat), .B(G203GAT_82_ngat), .Y(Ginternal__51gat) );
AND2XL U_g52 (.A(G180GAT_56_ngat), .B(G203GAT_82_gat), .Y(Ginternal__52gat) );
AND2XL U_g53 (.A(G102GAT_31_gat), .B(G213GAT_83_gat), .Y(G259GAT_86_gat) );
OR2XL U_g54 (.A(Ginternal__56gat), .B(Ginternal__55gat), .Y(G247GAT_87_gat) );
AND2XL U_g55 (.A(G177GAT_59_gat), .B(G203GAT_82_ngat), .Y(Ginternal__55gat) );
AND2XL U_g56 (.A(G177GAT_59_ngat), .B(G203GAT_82_gat), .Y(Ginternal__56gat) );
AND2XL U_g57 (.A(G89GAT_27_gat), .B(G213GAT_83_gat), .Y(G258GAT_88_gat) );
OR2XL U_g58 (.A(Ginternal__60gat), .B(Ginternal__59gat), .Y(G243GAT_89_gat) );
AND2XL U_g59 (.A(G174GAT_62_gat), .B(G203GAT_82_ngat), .Y(Ginternal__59gat) );
AND2XL U_g60 (.A(G174GAT_62_ngat), .B(G203GAT_82_gat), .Y(Ginternal__60gat) );
AND2XL U_g61 (.A(G76GAT_23_gat), .B(G213GAT_83_gat), .Y(G257GAT_90_gat) );
OR2XL U_g62 (.A(Ginternal__64gat), .B(Ginternal__63gat), .Y(G239GAT_91_gat) );
AND2XL U_g63 (.A(G171GAT_65_gat), .B(G203GAT_82_ngat), .Y(Ginternal__63gat) );
AND2XL U_g64 (.A(G171GAT_65_ngat), .B(G203GAT_82_gat), .Y(Ginternal__64gat) );
AND2XL U_g65 (.A(G63GAT_19_gat), .B(G213GAT_83_gat), .Y(G256GAT_92_gat) );
OR2XL U_g66 (.A(Ginternal__68gat), .B(Ginternal__67gat), .Y(G236GAT_93_gat) );
AND2XL U_g67 (.A(G168GAT_68_gat), .B(G203GAT_82_ngat), .Y(Ginternal__67gat) );
AND2XL U_g68 (.A(G168GAT_68_ngat), .B(G203GAT_82_gat), .Y(Ginternal__68gat) );
AND2XL U_g69 (.A(G50GAT_15_gat), .B(G213GAT_83_gat), .Y(G255GAT_94_gat) );
OR2XL U_g70 (.A(Ginternal__72gat), .B(Ginternal__71gat), .Y(G233GAT_95_gat) );
AND2XL U_g71 (.A(G165GAT_71_gat), .B(G203GAT_82_ngat), .Y(Ginternal__71gat) );
AND2XL U_g72 (.A(G165GAT_71_ngat), .B(G203GAT_82_gat), .Y(Ginternal__72gat) );
AND2XL U_g73 (.A(G37GAT_11_gat), .B(G213GAT_83_gat), .Y(G254GAT_96_gat) );
OR2XL U_g74 (.A(Ginternal__76gat), .B(Ginternal__75gat), .Y(G230GAT_97_gat) );
AND2XL U_g75 (.A(G162GAT_74_gat), .B(G203GAT_82_ngat), .Y(Ginternal__75gat) );
AND2XL U_g76 (.A(G162GAT_74_ngat), .B(G203GAT_82_gat), .Y(Ginternal__76gat) );
AND2XL U_g77 (.A(G24GAT_7_gat), .B(G213GAT_83_gat), .Y(G250GAT_98_gat) );
OR2XL U_g78 (.A(Ginternal__80gat), .B(Ginternal__79gat), .Y(G227GAT_99_gat) );
AND2XL U_g79 (.A(G159GAT_77_gat), .B(G203GAT_82_ngat), .Y(Ginternal__79gat) );
AND2XL U_g80 (.A(G159GAT_77_ngat), .B(G203GAT_82_gat), .Y(Ginternal__80gat) );
AND2XL U_g81 (.A(G11GAT_3_gat), .B(G213GAT_83_gat), .Y(G246GAT_100_gat) );
OR2XL U_g82 (.A(Ginternal__84gat), .B(Ginternal__83gat), .Y(G224GAT_101_gat) );
AND2XL U_g83 (.A(G154GAT_80_gat), .B(G203GAT_82_ngat), .Y(Ginternal__83gat) );
AND2XL U_g84 (.A(G154GAT_80_ngat), .B(G203GAT_82_gat), .Y(Ginternal__84gat) );
AND2XL U_g85 (.A(G213GAT_83_gat), .B(G1GAT_0_gat), .Y(G242GAT_102_gat) );
AND2XL U_g86 (.A(G198GAT_54_gat), .B(G251GAT_85_gat), .Y(G295GAT_103_gat) );
AND2XL U_g87 (.A(G197GAT_55_gat), .B(G251GAT_85_gat), .Y(G285GAT_104_gat) );
AND2XL U_g88 (.A(G196GAT_57_gat), .B(G247GAT_87_gat), .Y(G294GAT_105_gat) );
AND2XL U_g89 (.A(G195GAT_58_gat), .B(G247GAT_87_gat), .Y(G282GAT_106_gat) );
AND2XL U_g90 (.A(G194GAT_60_gat), .B(G243GAT_89_gat), .Y(G293GAT_107_gat) );
AND2XL U_g91 (.A(G193GAT_61_gat), .B(G243GAT_89_gat), .Y(G279GAT_108_gat) );
AND2XL U_g92 (.A(G192GAT_63_gat), .B(G239GAT_91_gat), .Y(G292GAT_109_gat) );
AND2XL U_g93 (.A(G191GAT_64_gat), .B(G239GAT_91_gat), .Y(G276GAT_110_gat) );
AND2XL U_g94 (.A(G190GAT_66_gat), .B(G236GAT_93_gat), .Y(G291GAT_111_gat) );
AND2XL U_g95 (.A(G189GAT_67_gat), .B(G236GAT_93_gat), .Y(G273GAT_112_gat) );
AND2XL U_g96 (.A(G188GAT_69_gat), .B(G233GAT_95_gat), .Y(G290GAT_113_gat) );
AND2XL U_g97 (.A(G187GAT_70_gat), .B(G233GAT_95_gat), .Y(G270GAT_114_gat) );
AND2XL U_g98 (.A(G186GAT_72_gat), .B(G230GAT_97_gat), .Y(G289GAT_115_gat) );
AND2XL U_g99 (.A(G185GAT_73_gat), .B(G230GAT_97_gat), .Y(G267GAT_116_gat) );
AND2XL U_g100 (.A(G184GAT_75_gat), .B(G227GAT_99_gat), .Y(G288GAT_117_gat) );
AND2XL U_g101 (.A(G183GAT_76_gat), .B(G227GAT_99_gat), .Y(G264GAT_118_gat) );
AND2XL U_g102 (.A(G158GAT_78_gat), .B(G224GAT_101_gat), .Y(G263GAT_119_gat) );
AND2XL U_g103 (.A(G157GAT_79_gat), .B(G224GAT_101_gat), .Y(G260GAT_120_gat) );
BUFX20 U_g104 (.A(G295GAT_103_gat), .Y(G308GAT_121_gat) );
AND9XL U_g105 (.A(G285GAT_104_gat), .B(G282GAT_106_gat), .C(G279GAT_108_gat), .D(G276GAT_110_gat), .E(G273GAT_112_gat), .F(G270GAT_114_gat), .G(G267GAT_116_gat), .H(G264GAT_118_gat), .I(G260GAT_120_gat), .Y(G296GAT_122_gat) );
BUFX20 U_g106 (.A(G294GAT_105_gat), .Y(G307GAT_123_gat) );
BUFX20 U_g107 (.A(G293GAT_107_gat), .Y(G306GAT_124_gat) );
BUFX20 U_g108 (.A(G292GAT_109_gat), .Y(G305GAT_125_gat) );
BUFX20 U_g109 (.A(G291GAT_111_gat), .Y(G304GAT_126_gat) );
BUFX20 U_g110 (.A(G290GAT_113_gat), .Y(G303GAT_127_gat) );
BUFX20 U_g111 (.A(G289GAT_115_gat), .Y(G302GAT_128_gat) );
BUFX20 U_g112 (.A(G288GAT_117_gat), .Y(G301GAT_129_gat) );
BUFX20 U_g113 (.A(G263GAT_119_gat), .Y(G300GAT_130_gat) );
BUFX20 U_g114 (.A(G296GAT_122_gat), .Y(G309GAT_131_gat) );
BUFX20 U_g115 (.A(G296GAT_122_gat), .Y(G319GAT_132_gat) );
BUFX20 U_g116 (.A(G296GAT_122_gat), .Y(G329GAT_133_gat) );
AND2XL U_g117 (.A(G112GAT_34_gat), .B(G319GAT_132_gat), .Y(G347GAT_134_gat) );
OR2XL U_g118 (.A(Ginternal__120gat), .B(Ginternal__119gat), .Y(G343GAT_135_gat) );
AND2XL U_g119 (.A(G285GAT_104_gat), .B(G309GAT_131_ngat), .Y(Ginternal__119gat) );
AND2XL U_g120 (.A(G285GAT_104_ngat), .B(G309GAT_131_gat), .Y(Ginternal__120gat) );
AND2XL U_g121 (.A(G99GAT_30_gat), .B(G319GAT_132_gat), .Y(G346GAT_136_gat) );
OR2XL U_g122 (.A(Ginternal__124gat), .B(Ginternal__123gat), .Y(G341GAT_137_gat) );
AND2XL U_g123 (.A(G282GAT_106_gat), .B(G309GAT_131_ngat), .Y(Ginternal__123gat) );
AND2XL U_g124 (.A(G282GAT_106_ngat), .B(G309GAT_131_gat), .Y(Ginternal__124gat) );
AND2XL U_g125 (.A(G86GAT_26_gat), .B(G319GAT_132_gat), .Y(G345GAT_138_gat) );
OR2XL U_g126 (.A(Ginternal__128gat), .B(Ginternal__127gat), .Y(G339GAT_139_gat) );
AND2XL U_g127 (.A(G279GAT_108_gat), .B(G309GAT_131_ngat), .Y(Ginternal__127gat) );
AND2XL U_g128 (.A(G279GAT_108_ngat), .B(G309GAT_131_gat), .Y(Ginternal__128gat) );
AND2XL U_g129 (.A(G73GAT_22_gat), .B(G319GAT_132_gat), .Y(G344GAT_140_gat) );
OR2XL U_g130 (.A(Ginternal__132gat), .B(Ginternal__131gat), .Y(G337GAT_141_gat) );
AND2XL U_g131 (.A(G276GAT_110_gat), .B(G309GAT_131_ngat), .Y(Ginternal__131gat) );
AND2XL U_g132 (.A(G276GAT_110_ngat), .B(G309GAT_131_gat), .Y(Ginternal__132gat) );
AND2XL U_g133 (.A(G60GAT_18_gat), .B(G319GAT_132_gat), .Y(G342GAT_142_gat) );
OR2XL U_g134 (.A(Ginternal__136gat), .B(Ginternal__135gat), .Y(G335GAT_143_gat) );
AND2XL U_g135 (.A(G273GAT_112_gat), .B(G309GAT_131_ngat), .Y(Ginternal__135gat) );
AND2XL U_g136 (.A(G273GAT_112_ngat), .B(G309GAT_131_gat), .Y(Ginternal__136gat) );
AND2XL U_g137 (.A(G47GAT_14_gat), .B(G319GAT_132_gat), .Y(G340GAT_144_gat) );
OR2XL U_g138 (.A(Ginternal__140gat), .B(Ginternal__139gat), .Y(G333GAT_145_gat) );
AND2XL U_g139 (.A(G270GAT_114_gat), .B(G309GAT_131_ngat), .Y(Ginternal__139gat) );
AND2XL U_g140 (.A(G270GAT_114_ngat), .B(G309GAT_131_gat), .Y(Ginternal__140gat) );
AND2XL U_g141 (.A(G34GAT_10_gat), .B(G319GAT_132_gat), .Y(G338GAT_146_gat) );
OR2XL U_g142 (.A(Ginternal__144gat), .B(Ginternal__143gat), .Y(G332GAT_147_gat) );
AND2XL U_g143 (.A(G267GAT_116_gat), .B(G309GAT_131_ngat), .Y(Ginternal__143gat) );
AND2XL U_g144 (.A(G267GAT_116_ngat), .B(G309GAT_131_gat), .Y(Ginternal__144gat) );
AND2XL U_g145 (.A(G21GAT_6_gat), .B(G319GAT_132_gat), .Y(G336GAT_148_gat) );
OR2XL U_g146 (.A(Ginternal__148gat), .B(Ginternal__147gat), .Y(G331GAT_149_gat) );
AND2XL U_g147 (.A(G264GAT_118_gat), .B(G309GAT_131_ngat), .Y(Ginternal__147gat) );
AND2XL U_g148 (.A(G264GAT_118_ngat), .B(G309GAT_131_gat), .Y(Ginternal__148gat) );
AND2XL U_g149 (.A(G319GAT_132_gat), .B(G8GAT_2_gat), .Y(G334GAT_150_gat) );
OR2XL U_g150 (.A(Ginternal__152gat), .B(Ginternal__151gat), .Y(G330GAT_151_gat) );
AND2XL U_g151 (.A(G260GAT_120_gat), .B(G309GAT_131_ngat), .Y(Ginternal__151gat) );
AND2XL U_g152 (.A(G260GAT_120_ngat), .B(G309GAT_131_gat), .Y(Ginternal__152gat) );
AND2XL U_g153 (.A(G308GAT_121_gat), .B(G343GAT_135_gat), .Y(G356GAT_152_gat) );
AND2XL U_g154 (.A(G307GAT_123_gat), .B(G341GAT_137_gat), .Y(G355GAT_153_gat) );
AND2XL U_g155 (.A(G306GAT_124_gat), .B(G339GAT_139_gat), .Y(G354GAT_154_gat) );
AND2XL U_g156 (.A(G305GAT_125_gat), .B(G337GAT_141_gat), .Y(G353GAT_155_gat) );
AND2XL U_g157 (.A(G304GAT_126_gat), .B(G335GAT_143_gat), .Y(G352GAT_156_gat) );
AND2XL U_g158 (.A(G303GAT_127_gat), .B(G333GAT_145_gat), .Y(G351GAT_157_gat) );
AND2XL U_g159 (.A(G302GAT_128_gat), .B(G332GAT_147_gat), .Y(G350GAT_158_gat) );
AND2XL U_g160 (.A(G301GAT_129_gat), .B(G331GAT_149_gat), .Y(G349GAT_159_gat) );
AND2XL U_g161 (.A(G300GAT_130_gat), .B(G330GAT_151_gat), .Y(G348GAT_160_gat) );
AND9XL U_g162 (.A(G356GAT_152_gat), .B(G355GAT_153_gat), .C(G354GAT_154_gat), .D(G353GAT_155_gat), .E(G352GAT_156_gat), .F(G351GAT_157_gat), .G(G350GAT_158_gat), .H(G349GAT_159_gat), .I(G348GAT_160_gat), .Y(G357GAT_161_gat) );
BUFX20 U_g163 (.A(G357GAT_161_gat), .Y(G360GAT_162_gat) );
BUFX20 U_g164 (.A(G357GAT_161_gat), .Y(G370GAT_163_gat) );
AND2XL U_g165 (.A(G115GAT_35_gat), .B(G360GAT_162_gat), .Y(G379GAT_164_gat) );
AND2XL U_g166 (.A(G105GAT_32_gat), .B(G360GAT_162_gat), .Y(G378GAT_165_gat) );
AND2XL U_g167 (.A(G92GAT_28_gat), .B(G360GAT_162_gat), .Y(G377GAT_166_gat) );
AND2XL U_g168 (.A(G79GAT_24_gat), .B(G360GAT_162_gat), .Y(G376GAT_167_gat) );
AND2XL U_g169 (.A(G66GAT_20_gat), .B(G360GAT_162_gat), .Y(G375GAT_168_gat) );
AND2XL U_g170 (.A(G53GAT_16_gat), .B(G360GAT_162_gat), .Y(G374GAT_169_gat) );
AND2XL U_g171 (.A(G40GAT_12_gat), .B(G360GAT_162_gat), .Y(G373GAT_170_gat) );
AND2XL U_g172 (.A(G27GAT_8_gat), .B(G360GAT_162_gat), .Y(G372GAT_171_gat) );
AND2XL U_g173 (.A(G360GAT_162_gat), .B(G14GAT_4_gat), .Y(G371GAT_172_gat) );
AND4XL U_g174 (.A(G108GAT_33_gat), .B(G379GAT_164_gat), .C(G347GAT_134_gat), .D(G259GAT_86_gat), .Y(G414GAT_173_gat) );
AND4XL U_g175 (.A(G95GAT_29_gat), .B(G378GAT_165_gat), .C(G346GAT_136_gat), .D(G258GAT_88_gat), .Y(G411GAT_174_gat) );
AND4XL U_g176 (.A(G82GAT_25_gat), .B(G377GAT_166_gat), .C(G345GAT_138_gat), .D(G257GAT_90_gat), .Y(G407GAT_175_gat) );
AND4XL U_g177 (.A(G69GAT_21_gat), .B(G376GAT_167_gat), .C(G344GAT_140_gat), .D(G256GAT_92_gat), .Y(G404GAT_176_gat) );
AND4XL U_g178 (.A(G56GAT_17_gat), .B(G375GAT_168_gat), .C(G342GAT_142_gat), .D(G255GAT_94_gat), .Y(G399GAT_177_gat) );
AND4XL U_g179 (.A(G43GAT_13_gat), .B(G374GAT_169_gat), .C(G340GAT_144_gat), .D(G254GAT_96_gat), .Y(G393GAT_178_gat) );
AND4XL U_g180 (.A(G30GAT_9_gat), .B(G373GAT_170_gat), .C(G338GAT_146_gat), .D(G250GAT_98_gat), .Y(G386GAT_179_gat) );
AND4XL U_g181 (.A(G17GAT_5_gat), .B(G372GAT_171_gat), .C(G336GAT_148_gat), .D(G246GAT_100_gat), .Y(G381GAT_180_gat) );
AND4XL U_g182 (.A(G371GAT_172_gat), .B(G334GAT_150_gat), .C(G242GAT_102_gat), .D(G4GAT_1_gat), .Y(G380GAT_181_gat) );
AND8XL U_g183 (.A(G414GAT_173_gat), .B(G411GAT_174_gat), .C(G407GAT_175_gat), .D(G404GAT_176_gat), .E(G399GAT_177_gat), .F(G393GAT_178_gat), .G(G386GAT_179_gat), .H(G381GAT_180_gat), .Y(G416GAT_182_gat) );
BUFX20 U_g184 (.A(G411GAT_174_gat), .Y(G420GAT_183_gat) );
BUFX20 U_g185 (.A(G407GAT_175_gat), .Y(G419GAT_184_gat) );
BUFX20 U_g186 (.A(G404GAT_176_gat), .Y(G418GAT_185_gat) );
BUFX20 U_g187 (.A(G393GAT_178_gat), .Y(G417GAT_186_gat) );
BUFX20 U_g188 (.A(G380GAT_181_gat), .Y(G415GAT_187_gat) );
AND2XL U_g189 (.A(G416GAT_182_ngat), .B(G415GAT_187_ngat), .Y(G421GAT_188_gat) );
AND4XL U_g190 (.A(G420GAT_183_gat), .B(G407GAT_175_gat), .C(G393GAT_178_gat), .D(G386GAT_179_gat), .Y(G429GAT_189_gat) );
AND4XL U_g191 (.A(G399GAT_177_gat), .B(G418GAT_185_gat), .C(G393GAT_178_gat), .D(G386GAT_179_gat), .Y(G425GAT_190_gat) );
AND3XL U_g192 (.A(G419GAT_184_gat), .B(G393GAT_178_gat), .C(G399GAT_177_gat), .Y(G428GAT_191_gat) );
AND2XL U_g193 (.A(G417GAT_186_gat), .B(G386GAT_179_gat), .Y(G422GAT_192_gat) );
AND4XL U_g194 (.A(G399GAT_177_gat), .B(G422GAT_192_gat), .C(G386GAT_179_gat), .D(G381GAT_180_gat), .Y(G430GAT_193_gat) );
AND4XL U_g195 (.A(G428GAT_191_gat), .B(G425GAT_190_gat), .C(G386GAT_179_gat), .D(G381GAT_180_gat), .Y(G431GAT_194_gat) );
AND4XL U_g196 (.A(G429GAT_189_gat), .B(G425GAT_190_gat), .C(G422GAT_192_gat), .D(G381GAT_180_gat), .Y(G432GAT_195_gat) );
INVXL U_g197 (.A(G115GAT_35_gat), .Y(G115GAT_35_ngat) );
INVXL U_g198 (.A(G151GAT_36_gat), .Y(G151GAT_36_ngat) );
INVXL U_g199 (.A(G112GAT_34_gat), .Y(G112GAT_34_ngat) );
INVXL U_g200 (.A(G105GAT_32_gat), .Y(G105GAT_32_ngat) );
INVXL U_g201 (.A(G147GAT_38_gat), .Y(G147GAT_38_ngat) );
INVXL U_g202 (.A(G99GAT_30_gat), .Y(G99GAT_30_ngat) );
INVXL U_g203 (.A(G92GAT_28_gat), .Y(G92GAT_28_ngat) );
INVXL U_g204 (.A(G143GAT_40_gat), .Y(G143GAT_40_ngat) );
INVXL U_g205 (.A(G86GAT_26_gat), .Y(G86GAT_26_ngat) );
INVXL U_g206 (.A(G79GAT_24_gat), .Y(G79GAT_24_ngat) );
INVXL U_g207 (.A(G139GAT_42_gat), .Y(G139GAT_42_ngat) );
INVXL U_g208 (.A(G73GAT_22_gat), .Y(G73GAT_22_ngat) );
INVXL U_g209 (.A(G66GAT_20_gat), .Y(G66GAT_20_ngat) );
INVXL U_g210 (.A(G135GAT_44_gat), .Y(G135GAT_44_ngat) );
INVXL U_g211 (.A(G60GAT_18_gat), .Y(G60GAT_18_ngat) );
INVXL U_g212 (.A(G53GAT_16_gat), .Y(G53GAT_16_ngat) );
INVXL U_g213 (.A(G131GAT_46_gat), .Y(G131GAT_46_ngat) );
INVXL U_g214 (.A(G47GAT_14_gat), .Y(G47GAT_14_ngat) );
INVXL U_g215 (.A(G40GAT_12_gat), .Y(G40GAT_12_ngat) );
INVXL U_g216 (.A(G127GAT_48_gat), .Y(G127GAT_48_ngat) );
INVXL U_g217 (.A(G34GAT_10_gat), .Y(G34GAT_10_ngat) );
INVXL U_g218 (.A(G27GAT_8_gat), .Y(G27GAT_8_ngat) );
INVXL U_g219 (.A(G123GAT_50_gat), .Y(G123GAT_50_ngat) );
INVXL U_g220 (.A(G21GAT_6_gat), .Y(G21GAT_6_ngat) );
INVXL U_g221 (.A(G14GAT_4_gat), .Y(G14GAT_4_ngat) );
INVXL U_g222 (.A(G119GAT_52_gat), .Y(G119GAT_52_ngat) );
INVXL U_g223 (.A(G8GAT_2_gat), .Y(G8GAT_2_ngat) );
INVXL U_g224 (.A(G203GAT_82_gat), .Y(G203GAT_82_ngat) );
INVXL U_g225 (.A(G180GAT_56_gat), .Y(G180GAT_56_ngat) );
INVXL U_g226 (.A(G177GAT_59_gat), .Y(G177GAT_59_ngat) );
INVXL U_g227 (.A(G174GAT_62_gat), .Y(G174GAT_62_ngat) );
INVXL U_g228 (.A(G171GAT_65_gat), .Y(G171GAT_65_ngat) );
INVXL U_g229 (.A(G168GAT_68_gat), .Y(G168GAT_68_ngat) );
INVXL U_g230 (.A(G165GAT_71_gat), .Y(G165GAT_71_ngat) );
INVXL U_g231 (.A(G162GAT_74_gat), .Y(G162GAT_74_ngat) );
INVXL U_g232 (.A(G159GAT_77_gat), .Y(G159GAT_77_ngat) );
INVXL U_g233 (.A(G154GAT_80_gat), .Y(G154GAT_80_ngat) );
INVXL U_g234 (.A(G309GAT_131_gat), .Y(G309GAT_131_ngat) );
INVXL U_g235 (.A(G285GAT_104_gat), .Y(G285GAT_104_ngat) );
INVXL U_g236 (.A(G282GAT_106_gat), .Y(G282GAT_106_ngat) );
INVXL U_g237 (.A(G279GAT_108_gat), .Y(G279GAT_108_ngat) );
INVXL U_g238 (.A(G276GAT_110_gat), .Y(G276GAT_110_ngat) );
INVXL U_g239 (.A(G273GAT_112_gat), .Y(G273GAT_112_ngat) );
INVXL U_g240 (.A(G270GAT_114_gat), .Y(G270GAT_114_ngat) );
INVXL U_g241 (.A(G267GAT_116_gat), .Y(G267GAT_116_ngat) );
INVXL U_g242 (.A(G264GAT_118_gat), .Y(G264GAT_118_ngat) );
INVXL U_g243 (.A(G260GAT_120_gat), .Y(G260GAT_120_ngat) );
INVXL U_g244 (.A(G415GAT_187_gat), .Y(G415GAT_187_ngat) );
INVXL U_g245 (.A(G416GAT_182_gat), .Y(G416GAT_182_ngat) );

endmodule
